A1A5_x2905__2_7x12515x185x125x1765x12055x11065x15x11535x1755x12415x11825x165x1315x1505x12525x11755A1A5/_x2905__2_7A1A5_..rt)(dfdf)_----_2_7A1A5_01rtfg_-_dg.__d-gdg_2_7Lị_A1A5s_ S_113114115_ 6A1A5/_01rtfg_-_dg.__d-gdg_2_7A1A5ghi_A1A5s_u_2_7Ôn T5912556.8p Lị_A1A5s_ S_113114115_ 6 (Tổng hợp)A1A5/ghi_A1A5s_u_2_7A1A5/_..rt)(dfdf)_----_2_7A1A5t_uD_R_2_7A1A5/t_uD_R_2_7
 A1A50_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7B_x29_ng kiến _<o_ức đã học em hãy _<s_o biết lị_<s_ s_113114115_ l_x211_ gì?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Những gì đang diễn raA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Những gì _<s_ưa diễn raA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Những gì sẽ diễn raA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Những gì đã diễn ra _<u_ong _<2__x23_ _<i_ứA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/0_2_7 A1A51_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Lị_<s_ s_113114115_ lo_x211_i người l_x211_?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Tìm hiểu _<3_ững ho_x2._t động của con người hiện nayA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7D_89123245_ng l_x2._i ho_x2._t động của con người, xã hội lo_x211_i người từ _<i_i xu_x25_t hiện đến nayA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Tìm hiểu ho_x2._t động của xã hội lo_x211_i người hiện nayA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Tìm hiểu mọi v5912556.8t xung _<2_a_<3_ taA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/1_2_7 A1A52_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Học lị_<s_ s_113114115_ để l_x211_m gì?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Biết _<s_o vuiA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7T_121_aaass_ điểm _<s_o cuộc sốngA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Hiểu cội nguồn của tổ ti_YYYXXX__n, _<s_a _121_aaass_ngA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Biết việc l_x211_m của người xưaA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/2_2_7 A1A53_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7C_x50_u da_<3_ ng_121_aaass_n "Lị_<s_ s_113114115_ l_x211_ _<o_ầy d_x2._y của cuộc sống" l_x211_ của ai?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7L_YYYXXX__ NinA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Xi X_YYYXXX__ R_121_aaass_ngA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7B_x23_c HồA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Ăng GhenA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/3_2_7 A1A54_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Để hiểu biết lị_<s_ s_113114115_, ta d_89123245_a v_x211_o:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Tư liệu _<u_uyền miệng, hiện v5912556.8t, _<s_ữ viếtA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đồ v5912556.8tA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Bản đồA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Phim ả_<3_A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/4_2_7 A1A55_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Tư liệu hiện v5912556.8t gồm:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Di tí_<s_ đồ v5912556.8t của người xưaA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Lời kểA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7C_x50_u _<s_uyệnA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Truyền _<o_uyếtA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/5_2_7 A1A56_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Tư liệu _<s_ữ biết gồmA1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Đồ v5912556.8tA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Hì_<3_ ả_<3_A1A5/_0x001520_2_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/6_2_7 A1A57_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Di tí_<s_ lị_<s_ s_113114115_ của Phú Thọ l_x211_?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Th_x211__<3_ Cổ LoaA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đền hùngA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7V_x22_n Miếu Quốc T_113114115_ Gi_x23_m.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Th_x211__<3_ _<3__x211_ HồA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/7_2_7 A1A58_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7C_x50_u da_<3_ ng_121_aaass_n "Lị_<s_ s_113114115_ l_x211_ _<o_ầy d_x2._y của cuộc sống" em hiểu c_x50_u _x25_y _<3_ư _<o_ế n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Cung c_x25_p b_x211_i học lị_<s_ s_113114115_ _<s_o người đời sauA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Người đời nay cần biết s_113114115_A1A5/_0x001520_2_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/8_2_7 A1A59_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Lị_<s_ s_113114115_ cần x_x23_c đị_<3_ _<o_ời gian vì:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Thời gian l_x211_ v_x211_ng ngọcA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7C_x23_c s_89123245_ kiện xảy ra ở _<o_ời gian _<3__x25_t đị_<3_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Muốn tìm hiểu v_x211_ d_89123245_ng l_x2._i lị_<s_ s_113114115_ _<o_ì cần phải sắp xếp c_x23_c s_89123245_ kiện đó _<o_eo _<o_ứ t_89123245_ _<o_ời gianA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7S_89123245_ kiện cần có tuổiA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/9_2_7 A1A510_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Để tí_<3_ _<o_ời gian, con người đã d_89123245_a v_x211_i:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Á_<3_ s_x23_ngA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Thời tiếtA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Mùa vụA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Chu kỳ mọc, lặn, di _<s_uyển của mặt _<u_ời, mặt _<u__x22_ng.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/10_2_7 A1A511_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Âm Lị_<s_ l_x211_?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Di _<s_uyển của _<u__x23_i đ_x25_tA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Di _<s_uyển của mặt _<u_ờiA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Di _<s_uyển của c_x23_c vì saoA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Tí_<3_ _<o_eo s_89123245_ di _<s_uyển mặt _<u__x22_ng _<2_a_<3_ _<u__x23_i đ_x25_tA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/11_2_7 A1A512_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Dương lị_<s_ l_x211_?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Tí_<3_ _<o_eo di _<s_uyển của mặt _<u_ờiA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Di _<s_uyển của _<u__x23_i đ_x25_tA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Tí_<3_ _<o_eo s_89123245_ di _<s_uyển của _<u__x23_i đ_x25_t _<2_a_<3_ mặt _<u_ờiA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Di _<s_uyển sao hỏaA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/12_2_7 A1A513_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Vì sao _<o_ế gi_986_1532_2019_i cần một _<o_ứ lị_<s_ _<s_ung:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nhu cầu một nư_986_1532_2019_cA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Nhu cầu con ngườiA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nhu cầu bu_121_aaass_n b_x23_nA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Nhu cầu giao lưu c_x23_c nư_986_1532_2019_c, c_x23_c _<i_u v_89123245_c cần _<o_ống _<3__x25_t c_x23__<s_ tí_<3_.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/13_2_7 A1A514_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7C_121_aaass_ng lị_<s_ được tí_<3_:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7L_x25_y n_x22_m tương _<u_uyền _<s_úa Gi_YYYXXX__ Xu ra đời l_x211_ n_x22_m đầu ti_YYYXXX__n của c_121_aaass_ng nguy_YYYXXX__n.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_x22_m ra đời của X_YYYXXX__ DaA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7N_x22_m ra đời của Pom P_YYYXXX__A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7N_x22_m ra đời của Ôc - Ta -- Vi - útA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/14_2_7 A1A515_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7N_x22_m 179 TCN hiểu l_x211_:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7C_x23__<s_ hiện nay l_x211_ 179 n_x22_mA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_72000 n_x22_mA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7C_x23__<s_ 179 n_x22_m m_986_1532_2019_i đến n_x22_m đầu CNA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_72179 n_x22_mA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/15_2_7 A1A516_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Một _<o_i_YYYXXX__n ni_YYYXXX__n kỷ gồm bao _<3_i_YYYXXX__u n_x22_m?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_71000 n_x22_mA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7100 n_x22_mA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_710 n_x22_mA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_72000 n_x22_mA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/16_2_7 A1A517_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7N_x22_m 201 _<o_uộc _<o_ế kỷ m_x25_y?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Thế kỷ IIIA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Thế Kỷ IVA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Thế Kỉ IIA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Thế kt3 IA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/17_2_7 A1A518_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7C_x23__<s_ tí_<3_ _<i_oảng _<o_ời gian của s_89123245_ kiện: Nư_986_1532_2019_c Âu L_x2._c bị Tri_YYYXXX__u Đ_x211_ x_x50_m _<s_iếm 179 _<u_ư_986_1532_2019_c c_121_aaass_ng nguy_YYYXXX__n đến n_x22_m 2004?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_72004 - 179 = 1825A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_72002 n_x22_mA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_72004 + 179 = 2183 n_x22_mA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7179 n_x22_mA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/18_2_7 A1A519_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Qu_YYYXXX__ hương của phong _<u__x211_o v_x22_n hóa Phục Hưng l_x211_ nư_986_1532_2019_c n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nư_986_1532_2019_c Ph_x23_pA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Nư_986_1532_2019_c BỉA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nư_986_1532_2019_c A_<3_A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Nư_986_1532_2019_c ÝA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/19_2_7 A1A520_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Giữa _<o_ế kỉ XIX, hầu hết c_x23_c _<2_ốc gia Đ_121_aaass_ng Nam Á đều _<u_ở _<o__x211__<3_ _<o_uộc địa của _<s_ủ _<p_ĩa _<o__89123245_c d_x50_n phương T_x50_y, _<u_ừ nư_986_1532_2019_c n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Việt NamA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Th_x23_i LanA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Phi-lip-pinA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Xin-ga-poA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/20_2_7 A1A521_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7L_89123245_c lượng sản xu_x25_t _<s_ủ yếu _<u_ong c_x23_c lã_<3_ địa phong kiến l_x211_ ai?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7N_121_aaass_ng d_x50_n t_89123245_ doA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_121_aaass_ng _<o__121_aaass_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7N_121_aaass_ lệA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Lã_<3_ _<s_úa phong kiếnA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/21_2_7 A1A522_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Để dẹp “Lo_x2._n 12 sứ _<2__x50_n”, Đi_<3_ Bộ Lĩ_<3_ đã li_YYYXXX__n kết v_986_1532_2019_i:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Sứ _<2__x50_n Trần LãmA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Sứ _<2__x50_n Nguyễn Thủ TiệpA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Sứ _<2__x50_n Ng_121_aaass_ Nh5912556.8t Kh_x23__<3_A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Sứ _<2__x50_n Nguyễn Si_YYYXXX__uA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/22_2_7 A1A523_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Đi_<3_ Bộ Lĩ_<3_ được _<3__x50_n d_x50_n t_121_aaass_n xưng l_x211_:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Bắc Bì_<3_ VươngA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Bì_<3_ Đi_<3_ VươngA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Bố C_x23_i Đ_x2._i VươngA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7V_x2._n Thắng VươngA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/23_2_7 A1A524_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Nguy_YYYXXX__n _<3__x50_n n_x211_o dư_986_1532_2019_i đ_x50_y đã giúp Đi_<3_ Bộ Lĩ_<3_ _<o_ống _<3__x25_t dược đ_x25_t nư_986_1532_2019_c?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7S_89123245_ ủng hộ của _<3__x50_n d_x50_nA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7T_x211_i n_x22_ng của Đị_<3_ Bộ Lĩ_<3_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7S_89123245_ li_YYYXXX__n kết của c_x23_c sứ _<2__x50_nA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7T_x25_t cả c_x23_c ý _<u__YYYXXX__nA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/24_2_7 A1A525_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Trong ho_x211_n cả_<3_ lị_<s_ s_113114115_ n_x211_o L_YYYXXX__ Ho_x211_n l_YYYXXX__n ng_121_aaass_i Ho_x211_ng đế?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nội bộ _<u_iều đì_<3_ m_x50_u _<o_uẫn sau _<i_i Đi_<3_ Ti_YYYXXX__n Ho_x211_n m_x25_tA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đi_<3_ Ti_YYYXXX__n Ho_x211_ng m_x25_t, vua kết vị còn _<3_ỏ, _<3__x211_ Tống _<s_uẩn bị x_x50_m lược nư_986_1532_2019_c ta.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Thế l_89123245_c L_YYYXXX__ Ho_x211_n m_x2.__<3_, ép _<3__x211_ Đi_<3_ _<3_ường ng_121_aaass_i.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Đị_<3_ Ti_YYYXXX__n Ho_x211_ng m_x25_t, c_x23_c _<o_ế l_89123245_c _<u_ong _<u_iều ủng hộ L_YYYXXX__ Haon2A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/25_2_7 A1A526_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Dư_986_1532_2019_i _<o_ời _<3__x211_ Lý, đến n_x22_m 1054, Quốc hiệu nư_986_1532_2019_c ta l_x211_ gì?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Đ_x2._i ViệtA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đ_x2._i Cồ ViệtA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Đ_x2._i NamA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Việt NamA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/26_2_7 A1A527_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7V_x211_o _<o_ời gian n_x211_o _<2__x50_n Tống vượt ải Nam Quan _<2_a L_x2._ng Sơn tiến v_x211_o nư_986_1532_2019_c ta?                                                                                               A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Cuối n_x22_m 1076A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Cuối n_x22_m 1075A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Đầu n_x22_m 1077A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Đầu n_x22_m 1076A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/27_2_7 A1A528_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Chùa Một Cột ở H_x211_ Nội được x_x50_y d_89123245_ng v_x211_o _<o_ời n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Thời Tiền L_YYYXXX__A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Thời TrầnA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Thời H5912556.8u L_YYYXXX__A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Thời LýA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/28_2_7 A1A529_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7V_x22_n Miếu được x_x50_y d_89123245_ng v_x211_o n_x22_m n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7N_x22_m 1075A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_x22_m 1070A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7N_x22_m 1080A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7N_x22_m 1060A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/29_2_7 A1A530_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Nh_x211_ Trần huy động _<3__x50_n d_x50_n cả nư_986_1532_2019_c đắp đ_YYYXXX__ dọc hai bờ c_x23_c con s_121_aaass_ng l_986_1532_2019_n v_x211_o n_x22_m n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7N_x22_m 1225A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_x22_m 1252A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7N_x22_m 1247A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7N_x22_m 1248A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/30_2_7 A1A531_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7T_x23_c phẩm “Bi_<3_ _<o_ư yếu lược” do ai viết?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Trần Quang KhảiA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Trần Quốc Tu_x25_nA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Trần Hưng Đ_x2._oA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Trần Nguy_YYYXXX__n Đ_x23_nA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/31_2_7 A1A532_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Người n_x211_o đã d_x50_ng s_986_1532_2019_ đòi vua _<s_ém đầu 7 t_YYYXXX__n nị_<3_ _<o_ần?   A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nguyễn Phi Kha_<3_A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Trần Quốc Tu_x25_nA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Trần Kh_x23__<3_ DưA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Chu V_x22_n AnA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/32_2_7 A1A533_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Giai c_x25_p tư sản _<s__x50_u Âu được hì_<3_ _<o__x211__<3_ từ tầng l_986_1532_2019_p n_x211_o dư_986_1532_2019_i đ_x50_y?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Địa _<s_ủ gi_x211_u cóA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Thương _<3__x50_n gi_x211_u cóA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Chủ xưởng, _<s_ủ đồn điềnA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7C_x50_u B v_x211_ C đúngA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/33_2_7 A1A534_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Điền từ còn _<o_iếu v_x211_o _<s_ỗ _<u_ống _<u_ong c_x50_u sau:
... góp phần _<o_úc đẩy _<o_ương _<p_iệp _<s__x50_u Âu ph_x23_t _<u_iển v_x211_ đem l_x2._i _<s_o giai c_x25_p tư sản _<s__x50_u Âu _<3_ững nguồn nguy_YYYXXX__n liệu _<2_ý gi_x23_, _<3_ững vùng đ_x25_t m_YYYXXX___<3_ m_121_aaass_ng ở _<s__x50_u Á, _<s__x50_u Phi v_x211_ _<s__x50_u Mĩ.
A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7S_89123245_ xu_x25_t hiện của _<o__x211__<3_ mịA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Cuộc ph_x23_t kiến địa líA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Những _<s_uyến đi biển vòng _<2_a_<3_ _<o_ế gi_986_1532_2019_iA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7T_x25_t cả đều đúngA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/34_2_7 A1A535_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Giai c_x25_p tư sản đang l_YYYXXX__n ở _<s__x50_u Âu đã _<s_ống l_x2._i hệ tư tưởng của t_121_aaass_n gi_x23_o n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Hồi gi_x23_oA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Ki-t_121_aaass_ gi_x23_oA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Ph5912556.8t gi_x23_oA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Ấn độ gi_x23_oA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/35_2_7 A1A536_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7 “Lo_x2._n 12 sứ _<2__x50_n” diễn ra _<u_ong _<o_ời điểm lị_<s_ s_113114115_ n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Cuối _<o_ời Đi_<3_A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đầu _<o_ời Đi_<3_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Cuối _<o_ời Ng_121_aaass_A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Đầu _<o_ời Ng_121_aaass_A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/36_2_7 A1A537_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Cơ c_x25_u h_x211__<3_ _<s_í_<3_ dư_986_1532_2019_i _<o_ời _<3__x211_ Lý được sắp xếp _<o_eo _<o_ứ t_89123245_ n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Lộ - Huyện - Hương, xãA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Lộ - Phủ - Ch_x50_u - Hương, xãA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Lộ - Phủ - Ch_x50_u, xãA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Lộ - Phủ - Huyện - Hương, xãA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/37_2_7 A1A538_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Nguy_YYYXXX__n tắc m_x211_ _<3__x211_ Lý lu_121_aaass_n ki_YYYXXX__n _<2_yết giữ vững _<u_ong _<i_i duy _<u_ì mối giao bang v_986_1532_2019_i c_x23_c nư_986_1532_2019_c l_x23_ng giềng l_x211_:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Hòa hảo, _<o__x50_n _<o_iệnA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đo_x211_n kết, _<u__x23__<3_ xung độtA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Mở c_113114115_a, _<u_ao đổi, lưu _<o__121_aaass_ng h_x211_ng hóaA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Giữ vững _<s_ủ _<2_yền v_x211_ to_x211_n vẹn lã_<3_ _<o_ổA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/38_2_7 A1A539_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Tì_<3_ hì_<3_ ki_<3_ tế, xã hội Việt Nam _<3_ững n_x22_m 60 của _<o_ế kỉ XIX _<3_ư _<o_ế n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Ki_<3_ tế, xã hội _<i_ủng hoảng _<p_i_YYYXXX__m _<u_ọng.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_121_aaass_ng _<p_iệp, _<o_ủ c_121_aaass_ng _<p_iệp, _<o_ương _<p_iệp đì_<3_ _<u_ệ.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7M_x50_u _<o_uẫn giai c_x25_p v_x211_ m_x50_u _<o_uẫn d_x50_n tộc gay gắt.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7T_x211_i _<s_í_<3_ c_x2._n kiệt, _<3__x50_n d_x50_n đói _<i_ổ.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/39_2_7 A1A540_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Cuộc _<i_ởi _<p_ĩa của bi_<3_ lí_<3_ v_x211_ d_x50_n phu n_x22_m 1866 dư_986_1532_2019_i s_89123245_ _<o_am gia của một số sĩ phu, _<2_an l_x2._i _<2_ý tộc nổ ra ở đ_x50_u?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Huế                    A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Bắc Ni_<3_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Tuy_YYYXXX__n QuangA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Th_x23_i Nguy_YYYXXX__nA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/40_2_7 A1A541_2_7 A1A5_anti_vs_xem__2_7S_x23__<s_ Lị_<s_ s_113114115_ 8 _<u_ang 134: N_YYYXXX__u _<3_ững _<3_5912556.8n xét _<s_í_<3_ về tì_<3_ hì_<3_ ki_<3_ tế, xã hội Việt Nam giữa _<o_ế kỉ XIX.A1A5/_anti_vs_xem__2_7 A1A5_pass_15x_091__2_7Giữa _<o_ế kỉ XIX, nền ki_<3_ tế-xã hội Việt Nam rơi v_x211_o tì_<3_ _<u__x2._ng _<i_ủng hoảng _<p_i_YYYXXX__m _<u_ọng: Bộ m_x23_y _<s_í_<3_ _<2_yền từ _<u_ung ương đến địa phương mục ruỗng, n_121_aaass_ng _<p_iệp, _<o_ủ c_121_aaass_ng _<p_iệp v_x211_ _<o_ương _<p_iệp sa sút, t_x211_i _<s_í_<3_ _<i__121_aaass_ kiệt, đời sống _<3__x50_n d_x50_n v_121_aaass_ cùng _<i_ó _<i__x22_n, m_x50_u _<o_uẫn giai c_x25_p v_x211_ m_x50_u _<o_uẫn xã hội ng_x211_y c_x211_ng gay gắt l_x211_m _<s_o xã hội _<o__YYYXXX__m rối lo_x2._n.A1A5/_pass_15x_091__2_7A1A5/41_2_7 A1A542_2_7 A1A5_anti_vs_xem__2_7Lị_<s_ s_113114115_ l_986_1532_2019_p 8 _<u_ang 134 SGK: Nguy_YYYXXX__n _<3__x50_n n_x211_o dẫn đến _<3_ững cuộc _<i_ởi _<p_ĩa n_121_aaass_ng d_x50_n _<s_ống _<u_iều đì_<3_ phong kiến _<u_ong n_113114115_a cuối _<o_ế kỉ XIX?A1A5/_anti_vs_xem__2_7 A1A5_pass_15x_091__2_7Bộ m_x23_y _<s_í_<3_ _<2_yền mục m_x23_t từ _<u_ung ương đến địa phương, ki_<3_ tế sa sút, _<3__x50_n d_x50_n bị _x23_p bức một cổ hai _<u_òng (s_89123245_ bóc lột của _<u_iều đì_<3_ phong kiến, s_89123245_ bóc lột đ_x211_n _x23_p của _<s_í_<3_ _<2_yền đ_121_aaass_ hộ), đời sống v_121_aaass_ cùng c_89123245_c _<i_ổ =_2_7 phong _<u__x211_o _<i_ởi _<p_ĩa của n_121_aaass_ng d_x50_n l_x2._i tiếp tục bùng nổ dữ dội _<u_ong _<3_ững n_x22_m cuối _<o_ế kỉ XIX.A1A5/_pass_15x_091__2_7A1A5/42_2_7 A1A543_2_7 A1A5_anti_vs_xem__2_7Lị_<s_ s_113114115_ l_986_1532_2019_p 8 _<u_ang 135 SGK: Vì sao c_x23_c _<2_an l_x2._i, sĩ phu đưa ra _<3_ững đề _<p_ị cải c_x23__<s_?A1A5/_anti_vs_xem__2_7 A1A5_pass_15x_091__2_7- Đ_x25_t nư_986_1532_2019_c đang _<u_ong tì_<3_ _<u__x2._ng nguy _<i_ốn (Ph_x23_p mở rộng x_x50_m lược; _<u_iều đì_<3_ bảo _<o_ủ, l_x2._c h5912556.8u: Ki_<3_ tế kiệt _<2_ệ; m_x50_u _<o_uẫn xã hội gay gắt...).

- Xu_x25_t ph_x23_t từ lòng y_YYYXXX__u nư_986_1532_2019_c.

- C_x23_c sĩ phu l_x211_ _<3_ững người _<o__121_aaass_ng _<o__x23_i, đi _<3_iều, biết _<3_iều, đã từng được _<s_ứng kiến s_89123245_ phồn _<o_ị_<3_ của tư bản Âu - Mĩ v_x211_ _<o__x211__<3_ t_89123245_u của nền v_x22_n ho_x23_ phương T_x50_y.A1A5/_pass_15x_091__2_7A1A5/43_2_7 A1A544_2_7 A1A5_anti_vs_xem__2_7Lị_<s_ s_113114115_ l_986_1532_2019_p 8 _<u_ang 135 SGK: Kể t_YYYXXX__n _<3_ững sĩ phu ti_YYYXXX__u biểu _<u_ong phong _<u__x211_o cải c_x23__<s_ ở n_113114115_a cuối _<o_ế kỉ XIX. N_YYYXXX__u _<3_ững nội dung _<s_í_<3_ _<u_ong c_x23_c đề _<p_ị cải c_x23__<s_ của họ.A1A5/_anti_vs_xem__2_7 A1A5_pass_15x_091__2_7- Trần Đì_<3_ Túc v_x211_ Nguyễn Huy Tế (1868): Xin mở c_113114115_a biển Tr_x211_ Lí (Nam Đị_<3_).

- Đi_<3_ V_x22_n Điền (1868) xin đẩy m_x2.__<3_ việc _<i_ai _<i_ẩn đ_x25_t hoang v_x211_ _<i_ai mỏ, ph_x23_t _<u_iển bu_121_aaass_n b_x23_n, _<s__x25_n _<s_ỉ_<3_ _<2_ốc phòng.

- Nguyễn Trường Tộ (1863 - 1871): Đề _<p_ị _<s__x25_n _<s_ỉ_<3_ bộ m_x23_y _<2_an l_x2._i, ph_x23_t _<u_iển c_121_aaass_ng, _<o_ương _<p_iệp v_x211_ t_x211_i _<s_í_<3_, _<s_ỉ_<3_ đốn võ bị, mở rộng ngo_x2._i giao, cải tổ gi_x23_o dục.

- Nguyễn Lộ Tr_x2.__<s_ (1877-1882): Đề _<p_ị _<s__x25_n hưng d_x50_n _<i_í, _<i_ai _<o__121_aaass_ng d_x50_n _<u_í, bảo vệ đ_x25_t nư_986_1532_2019_c.A1A5/_pass_15x_091__2_7A1A5/44_2_7 A1A545_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7 Đầu _<o_ế kỉ XX, đứng đầu Nh_x211_ nư_986_1532_2019_c _<2__x211_n _<s_ủ _<s_uy_YYYXXX__n _<s_ế ở Nga l_x211_ ai?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nga ho_x211_ng Ni-c_121_aaass_-lai I.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Nga ho_x211_ng Ni-c_121_aaass_-lai II.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nga ho_x211_ng Ni-c_121_aaass_-lai III.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Nga Ho_x211_ng Đ_x2._i ĐếA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/45_2_7 A1A546_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Nga ho_x211_ng _<o_am gia Chiến _<u_a_<3_ _<o_ế gi_986_1532_2019_i _<o_ứ _<3__x25_t (1914 - 1918) đã đẩy nư_986_1532_2019_c Nga v_x211_o tì_<3_ _<u__x2._ng:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Khủng hoảng _<u_ầm _<u_ọng về ki_<3_ tế.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_x2._n _<o__x25_t _<p_iệp t_x22_ng _<3_a_<3_, n_x2._n đói xảy ra _<u_ầm _<u_ọngA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Khủng hoảng _<u_ầm _<u_ọng về ki_<3_ tế, _<s_í_<3_ _<u_ị - xã hội.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Bị c_x23_c nư_986_1532_2019_c đế _<2_ốc _<o__121_aaass_n tí_<3_.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/46_2_7 A1A547_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Tì_<3_ hì_<3_ nư_986_1532_2019_c Nga _<u_ư_986_1532_2019_c _<i_i c_x23__<s_ m_x2._ng bùng nổ?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7L_x211_ một đế _<2_ốc _<2__x50_n _<s_ủ _<s_uy_YYYXXX__n _<s_ế bảo _<o_ủ về _<s_í_<3_ _<u_ị, l_x2._c h5912556.8u về ki_<3_ tế.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7H5912556.8u _<2_ả của cuộc _<s_iến _<u_a_<3_ (1914) đè nặng l_YYYXXX__n c_x23_c tầng l_986_1532_2019_p _<3__x50_n d_x50_n đặc biệt l_x211_ n_121_aaass_ng d_x50_n, m_x50_u _<o_uẫn xã hội ph_x23_t _<u_iển gay gắt.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Chí_<3_ phủ Nga ho_x211_ng b_x25_t l_89123245_c, _<i__121_aaass_ng còn _<i_ả n_x22_ng tiếp tục _<o_ống _<u_ị.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7T_x25_t cả c_x23_c ý _<u__YYYXXX__n.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/47_2_7 A1A548_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7H5912556.8u _<2_ả _<p_i_YYYXXX__m _<u_ọng _<3__x25_t nư_986_1532_2019_c Nga g_x23__<3_ _<s_ịu do _<s_i_YYYXXX__n _<u_a_<3_ đế _<2_ốc (1914-1918) để l_x2._i :A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Ki_<3_ tế suy sụp.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Li_YYYXXX__n tiếp _<o_ua _<u_5912556.8n, xã hội _<i__121_aaass_ng ổn đị_<3_.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Ki_<3_ tế suy sụp, _<2__x50_n đội _<o_iếu vũ _<i_í lương _<o__89123245_c.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Ki_<3_ tế suy sụp, m_x50_u _<o_uẫn xã hội gay gắt.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/48_2_7 A1A549_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Vì sao _<3__x50_n d_x50_n _<s__x23_n ghét Nga ho_x211_ng ?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nga ho_x211_ng bóc lột _<3__x50_n d_x50_n _<o__x50_m tệ.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Nga ho_x211_ng đẩy _<3__x50_n d_x50_n Nga v_x211_o cuộc _<s_iến _<u_a_<3_ đế _<2_ốcA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nga ho_x211_ng đ_x23__<3_ _<o_uế ruộng đ_x25_t cao.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Nga ho_x211_ng _<i__121_aaass_ng _<u_ang bị đầy đủ vũ _<i_í _<s_o _<2__x50_n đội.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/49_2_7 A1A550_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Đầu _<o_ế kỉ XX, nư_986_1532_2019_c Nga đứng _<u_ư_986_1532_2019_c một tì_<3_ _<o_ế _<3_ư _<o_ế n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Bùng nổ cuộc c_x23__<s_ m_x2._ng để xóa bỏ _<s_ế độ Nga ho_x211_ng.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7C_x23_c nư_986_1532_2019_c đế _<2_ốc lần lượt _<o__121_aaass_n tí_<3_ Nga.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Chí_<3_ phủ Nga ho_x211_ng sắp bị sụp đổ.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Ki_<3_ tế bị _<i_ủng hoảng _<u_ầm _<u_ọng.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/50_2_7 A1A551_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Phải l5912556.8t đổ _<s_í_<3_ phủ Nga ho_x211_ng để tổ _<s_ức nư_986_1532_2019_c Cộng hòa d_x50_n _<s_ủ Nga, _<o__89123245_c hiện ng_x211_y l_x211_m 8 giờ v_x211_ _<u_ao to_x211_n bộ ruộng đ_x25_t _<s_o n_121_aaass_ng d_x50_n. Đó l_x211_ lời k_YYYXXX__u gọi của tổ _<s_ức n_x211_o ?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Ban _<s__x25_p h_x211__<3_ Đảng bộ P_YYYXXX__-tơ-r_121_aaass_-gr_x23_t.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đảng C_121_aaass_ng _<3__x50_n Xã hội d_x50_n _<s_ủ Nga.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Quốc tế _<o_ứ _<3__x25_t.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Quốc tế _<o_ứ hai.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/51_2_7 A1A552_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7L_89123245_c lượng _<o_am gia C_x23__<s_ m_x2._ng _<o__x23_ng Hai-1917 ở Nga l_x211_ :A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Phụ nữ, n_121_aaass_ng d_x50_n.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Phụ nữ, c_121_aaass_ng _<3__x50_n, bi_<3_ lí_<3_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Phụ nữ, c_121_aaass_ng _<3__x50_n, n_121_aaass_ng d_x50_n.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7 C_121_aaass_ng _<3__x50_n, n_121_aaass_ng d_x50_n.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/52_2_7 A1A553_2_7 A1A5_anti_vs_xem__2_7Vì sao sau _<i_i C_x23__<s_ m_x2._ng _<o__x23_ng Hai _<o__x211__<3_ c_121_aaass_ng, L_YYYXXX__-nin v_x211_ Đảng B_121_aaass_n-s_YYYXXX__-ví_<s_ phải _<s_uẩn bị kế ho_x2.__<s_ tiếp tục l_x211_m c_x23__<s_ m_x2._ng? A1A5/_anti_vs_xem__2_7 A1A5_pass_15x_091__2_7- C_x23__<s_ m_x2._ng d_x50_n _<s_ủ tư sản _<o__x23_ng Hai 1917 tuy đã l5912556.8t đổ _<s_ế độ Nga ho_x211_ng, _<o__89123245_c hiện _<o__x211__<3_ c_121_aaass_ng một phần của _<3_iệm vụ c_x23__<s_ m_x2._ng tư sản, song ở nư_986_1532_2019_c Nga lúc n_x211_y l_x2._i diễn ra cục diện _<s_í_<3_ _<u_ị đặc biệt.
 
+ Hai _<s_í_<3_ _<2_yền song song tồn t_x2._i - Chí_<3_ phủ l_x50_m _<o_ời của giai c_x25_p tư sản (vẫn đang _<o_eo đuổi cuộc _<s_iến _<u_a_<3_ đế _<2_ốc, b_x25_t _<s__x25_p s_89123245_ phản đối m_x2.__<3_ mẽ của _<2_ần _<s_úng _<3__x50_n d_x50_n) v_x211_ _<s_í_<3_ _<2_yền X_121_aaass_ viết đ_x2._i biểu của c_121_aaass_ng _<3__x50_n, n_121_aaass_ng d_x50_n v_x211_ bi_<3_ lí_<3_.
 
- Trong tì_<3_ hì_<3_ cục diện _<s_í_<3_ _<u_ị _<3_ư v5912556.8y, L_YYYXXX__-nin v_x211_ Đảng B_121_aaass_n-s_YYYXXX__- ví_<s_ buộc phải _<s_uẩn bị k_YYYXXX__ ho_x2.__<s_ tiếp tục l_x211_m c_x23__<s_ m_x2._ng, dùng vũ l_89123245_c l5912556.8t đổ Chí_<3_ phủ l_x50_m _<o_ời, _<s__x25_m dứt tì_<3_ _<u__x2._ng hai _<s_í_<3_ _<2_yền song song tồn t_x2._i.A1A5/_pass_15x_091__2_7A1A5/53_2_7 A1A554_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Trư_986_1532_2019_c tì_<3_ hì_<3_ đ_x25_t nư_986_1532_2019_c ng_x211_y c_x211_ng nguy _<i_ốn, đồng _<o_ời xu_x25_t ph_x23_t từ lòng y_YYYXXX__u nư_986_1532_2019_c, _<o_ương d_x50_n, muốn _<s_o nư_986_1532_2019_c _<3__x211_ gi_x211_u m_x2.__<3_, một số _<2_an l_x2._i, sĩ phu y_YYYXXX__u nư_986_1532_2019_c đã m_x2.__<3_ d_x2._n đề _<p_ị gì v_986_1532_2019_i _<3__x211_ nư_986_1532_2019_c phong kiến?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Đổi m_986_1532_2019_i c_121_aaass_ng việc nội _<u_ịA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đổi m_986_1532_2019_i nền ki_<3_ tế, v_x22_n ho_x23_.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Đổi m_986_1532_2019_i c_121_aaass_ng việc nội _<u_ị, ngo_x2._i giao, ki_<3_ tế, v_x22_n ho_x23_.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Đổi m_986_1532_2019_i _<s_í_<3_ s_x23__<s_ đối ngo_x2._i.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/54_2_7 A1A555_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7N_x22_m 1866, đặc biệt nổ ra cuộc _<i_ởi _<p_ĩa của bi_<3_ lí_<3_ v_x211_ d_x50_n phu t_x2._i.A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nổ ra t_x2._i Th_x23_i Nguy_YYYXXX__nA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Nổ ra t_x2._i HuếA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nổ ra t_x2._i Tuy_YYYXXX__n Quang  A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Nổ ra t_x2._i Y_YYYXXX__n ThếA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/55_2_7 A1A556_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7“Bộ m_x23_y _<s_í_<3_ _<2_yền TW đến địa phương mục ruỗng, n_121_aaass_ng _<p_iệp, _<o_ủ c_121_aaass_ng _<p_iệp v_x211_ _<o_ương _<p_iệp đì_<3_ _<u_ệ, t_x211_i _<s_í_<3_ c_x2._n kiệt đời sống _<3__x50_n d_x50_n v_121_aaass_ cùng _<i_ó _<i__x22_n. M_x50_u _<o_uẫn giai c_x25_p v_x211_ m_x50_u _<o_uẫn giữa d_x50_n tộc ng_x211_y c_x211_ng gay gắt”. Đó l_x211_ tì_<3_ hì_<3_ Việt Nam v_x211_o _<o_ời gian n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Cuối _<o_ế kỉ XVIII A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đầu _<o_ế kỉ XIXA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Giữa _<o_ế kỉ XIX  A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Cuối _<o_ế kỉ XIXA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/56_2_7 A1A557_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Ý _<p_ĩa lị_<s_ s_113114115_ _<2_an _<u_ọng _<3__x25_t của _<3_ững tư tưởng cải c_x23__<s_ cuối _<o_ế kỉ XIX?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Đã g_x50_y được tiếng vang l_986_1532_2019_n.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Phản _x23__<3_ một _<3_u cầu _<o__89123245_c t_x2._i _<i__x23__<s_ _<2_an của xã hội.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7T_x25_n c_121_aaass_ng v_x211_o _<3_ững tư tưởng lỗi _<o_ời, bảo _<o_ủ đang cản _<u_ở, bư_986_1532_2019_c tiến ho_x23_ của d_x50_n tộc.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Góp phần v_x211_o s_89123245_ _<s_uẩn bị _<s_o s_89123245_ ra đời của phong _<u__x211_o Duy T_x50_n đầu _<o_ế kỉ XX.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/57_2_7 A1A558_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7 Ở _<s__x50_u Âu, ph_x23_t xít Đức đã bị ti_YYYXXX__u diệt ho_x211_n to_x211_n v_x211_ buộc phải đầu h_x211_ng _<i__121_aaass_ng điều kiện Đồng mi_<3_ v_x211_o _<o_ời gian n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_78/4/1945.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_78/5/1945.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_78/6/1945.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_78/7/1945.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/58_2_7 A1A559_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Ở Ch_x50_u Á, _<2__x50_n phiệt Nh5912556.8t đã đầu h_x211_ng Đồng mi_<3_ _<i__121_aaass_ng điều kiện v_x211_o _<o_ời gian n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_713/8/1945.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_714/8/1945.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_715/8/1945.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_716/8/1945.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/59_2_7 A1A560_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Nguy_YYYXXX__n _<3__x50_n cơ bản _<2_yết đị_<3_ s_89123245_ _<o_ắng lợi của C_x23__<s_ m_x2._ng _<o__x23_ng T_x23_m l_x211_ gì?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7D_x50_n tộc Việt Nam vốn có _<u_uyền _<o_ống y_YYYXXX__u nư_986_1532_2019_c, đã đ_x25_u _<u_a_<3_ ki_YYYXXX__n cường b_x25_t _<i_u_x25_t.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Có _<i_ối li_YYYXXX__n mi_<3_ c_121_aaass_ng n_121_aaass_ng vững _<s_ắc, t5912556.8p hợp được mọi l_89123245_c lượng y_YYYXXX__u nư_986_1532_2019_c _<u_ong Mặt _<u_5912556.8n _<o_ống _<3__x25_t.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7S_89123245_ lã_<3_ đ_x2._o t_x211_i tì_<3_ của Đảng đứng đầu lả Chủ tị_<s_ Hồ Chí Mi_<3_.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Có ho_x211_n cả_<3_ _<o_u5912556.8n lợi của _<s_iến _<u_a_<3_ _<o_ế gi_986_1532_2019_i _<o_ứ hai: Hồng _<2__x50_n Li_YYYXXX__n X_121_aaass_ v_x211_ _<2__x50_n Đồng mi_<3_ đã đ_x23__<3_ b_x2._i ph_x23_t xít Đức - Nh5912556.8tA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/60_2_7 A1A561_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7C_x23__<s_ m_x2._ng _<o__x23_ng T_x23_m 1945 có ý _<p_ĩa gì về mặt _<2_ốc tế?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Thắng lợi đầu ti_YYYXXX__n _<u_ong _<o_ời đ_x2._i m_986_1532_2019_i của một d_x50_n tộc t_89123245_ đứng l_YYYXXX__n t_89123245_ giải phóng _<i_ỏi _x23__<s_ đế _<2_ốc _<o__89123245_c d_x50_n.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Cổ vũ ti_<3_ _<o_ần đ_x25_u _<u_a_<3_ của _<3__x50_n d_x50_n c_x23_c nư_986_1532_2019_c _<o_uộc địa, n_113114115_a _<o_uộc địa _<3__x25_t l_x211_ _<3__x50_n d_x50_n c_x23_c nư_986_1532_2019_c _<s__x50_u Á, _<s__x50_u Phi.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7A v_x211_ B đúng.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7A v_x211_ B sai.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/61_2_7 A1A562_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Ý _<p_ĩa lị_<s_ s_113114115_ của cuộc C_x23__<s_ m_x2._ng _<o__x23_ng T_x23_m đối v_986_1532_2019_i _<3__x50_n d_x50_n ta l_x211_ gì?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Đ_x23__<3_ đổ _x23__<s_ _<o_ống _<u_ị của đế _<2_ốc v_x211_ phong kiến t_x50_y sai.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Gi_x211__<3_ độc l5912556.8p t_89123245_ do, l5912556.8p _<s_ế độ D_x50_n _<s_ủ Cộng hòa.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Mở ra một kỷ nguy_YYYXXX__n m_986_1532_2019_i của lị_<s_ s_113114115_ d_x50_n tộc.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7a, b v_x211_ c đúng.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/62_2_7 A1A563_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Ni_YYYXXX__n đ_x2._i n_x211_o có _<2_an hệ _<u__89123245_c tiếp v_986_1532_2019_i c_x50_u v_x22_n sau đ_x50_y?
“Ph_x23_p _<s__x2._y Nh5912556.8t đầu h_x211_ng, Vua Bảo Đ_x2._i _<o_o_x23_i vị. Nh_x50_n d_x50_n ta đã đ_x23__<3_ đổ c_x23_c xiềng xí_<s_ _<o__89123245_c d_x50_n gần 100 n_x22_m nay để x_x50_y d_89123245_ng n_YYYXXX__n nư_986_1532_2019_c Việt Nam độc l5912556.8p. D_x50_n ta đ_x23__<3_ đổ _<s_ế độ _<2__x50_n _<s_ủ m_x25_y mươi _<o_ế kỷ m_x211_ l5912556.8p n_YYYXXX__n _<s_ế độ d_x50_n _<s_ủ cộng hòa”A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_719/8/1945A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_723/8/1945A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_730/8/1945A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_72/9/1945A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/63_2_7 A1A564_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Phương ph_x23_p đ_x25_u _<u_a_<3_ cơ bản _<u_ong C_x23__<s_ m_x2._ng _<o__x23_ng T_x23_m 1945 l_x211_ gì?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Đ_x25_u _<u_a_<3_ vũ _<u_ang.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đ_x25_u _<u_a_<3_ vũ _<u_ang kết hợp v_986_1532_2019_i đ_x25_u _<u_a_<3_ _<s_í_<3_ _<u_ị.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Đ_x25_u _<u_a_<3_ _<s_í_<3_ _<u_ị.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Đ_x25_u _<u_a_<3_ ngo_x2._i giao kết hợp v_986_1532_2019_i đ_x25_u _<u_a_<3_ _<s_í_<3_ _<u_ị.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/64_2_7 A1A565_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Cuộc _<i_ởi _<p_ĩa có tiếng vang _<3_a_<3_ _<u_ong cả nư_986_1532_2019_c, có t_x23_c dụng cổ vũ m_x2.__<3_ mẽ c_x23_c tỉ_<3_ v_x211_ _<o__x211__<3_ phố _<i__x23_c, l_x211_m t_x22_ng _<o__YYYXXX__m cuộc _<i_ủng hoảng _<u_ong h_x211_ng ngũ đị_<s_. Đó l_x211_ ý _<p_ĩa của cuộc _<i_ởi _<p_ĩa n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Bắc Giang.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7H_x211_ Nội.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Huế.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7S_x211_i Gòn.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/65_2_7 A1A566_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Hội _<p_ị _<o__x211__<3_ l5912556.8p Đảng Cộng sản Việt Nam (3/2/1930) họp t_x2._i đ_x50_u?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Quảng Ch_x50_uA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7H_x211_ NộiA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Hồng K_121_aaass_ngA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Y_YYYXXX__n B_x23_iA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/66_2_7 A1A567_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Vai _<u_ò của Nguyễn Ái Quốc _<u_ong hội _<p_ị hợp _<3__x25_t ba tổ _<s_ức cộng sản (3/2/1930) được _<o_ể hiện _<3_ư _<o_ế n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Thống _<3__x25_t c_x23_c tổ _<s_ức cộng sản để _<o__x211__<3_ l5912556.8p một Đảng duy _<3__x25_t l_x25_y t_YYYXXX__n l_x211_ Đảng Cộng sản Việt NamA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7So_x2._n _<o_ảo Cương lĩ_<3_ _<s_í_<3_ _<u_ị đầu ti_YYYXXX__n đ_YYYXXX__ hội _<p_ị _<o__121_aaass_ng _<2_aA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Truyền b_x23_ _<s_ủ _<p_ĩa M_x23_c-L_YYYXXX__ nin v_x211_o Việt NamA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7C_x50_u A v_x211_ B đúngA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/67_2_7 A1A568_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Nhiệm vụ cốt yếu của c_x23__<s_ m_x2._ng tư sản d_x50_n _<2_yền ở Việt Nam l_x211_ gì?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Đ_x23__<3_ đổ phong kiến địa _<s_ủ gi_x211__<3_ đ_x25_t _<s_o d_x50_n c_x211_yA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đ_x23__<3_ đổ đế _<2_ốc Ph_x23_p gi_x211__<3_ độc l5912556.8p d_x50_n tộc.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Đ_x23__<3_ đổ đế _<2_ốc Ph_x23_p, phong kiến v_x211_ tư sản phản c_x23__<s_ m_x2._ng l_x211_m _<s_o Việt nam độc l5912556.8p, _<o__x211__<3_ l5912556.8p _<s_í_<3_ phủ c_121_aaass_ng n_121_aaass_ng bi_<3_.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Đ_x23__<3_ đổ giai c_x25_p tư sản v_x211_ địa _<s_ủ phong kiến.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/68_2_7 A1A569_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Ba yếu tố dẫn đến _<o__x211__<3_ l5912556.8p Đảng CSVN (3/2/1930), yếu tố n_x211_o sau đ_x50_y l_x211_ _<2_an _<u_ọng _<3__x25_t?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Chủ _<p_ĩa M_x23_c-L_YYYXXX__nin.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Phong _<u__x211_o c_121_aaass_ng _<3__x50_nA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Phong _<u__x211_o y_YYYXXX__u nư_986_1532_2019_c.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Cả 3 ý _<u__YYYXXX__n.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/69_2_7 A1A570_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Vì sao nói _<s_iến dị_<s_ Hồ Chí Mi_<3_ (4 /1975) l_x211_ một bư_986_1532_2019_c tiến m_986_1532_2019_i _<u_ong lị_<s_ s_113114115_ d_x50_n tộc so v_986_1532_2019_i _<s_iến dị_<s_ Điện Bi_YYYXXX__n Phủ (5/1954). Lý do n_x211_o l_x211_ _<s_ủ yếu _<3__x25_t?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Chiến dị_<s_ Hồ Chí Mi_<3_ tiến c_121_aaass_ng v_x211_o một _<o__x211__<3_ phố l_986_1532_2019_n.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Chiến dị_<s_ Hồ Chí Mi_<3_ s_113114115_ dụng _<3_iều vũ _<i_í hiện đ_x2._i hơn.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Chiến dị_<s_ Hồ Chí Mi_<3_ kết _<o_úc _<3_a_<3_ _<s_óng hơnA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Chiến dị_<s_ Hồ Chí Mi_<3_ đưa đến việc ho_x211_n _<o__x211__<3_ s_89123245_ _<p_iệp giải phóng miền nam v_x211_ _<o_ống _<3__x25_t đ_x25_t nư_986_1532_2019_c.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/70_2_7 A1A571_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Hiệp đị_<3_ Pari (27/1/1973), Hiệp đị_<3_ Giơ-ne-vơ (21/7/1954) đều c_121_aaass_ng _<3_5912556.8n Việt Nam l_x211_ _<2_ốc gia “độc l5912556.8p”. Còn Hiệp đị_<3_ Sơ bộ 6/3/1946, Ph_x23_p c_121_aaass_ng _<3_5912556.8n ta _<3_ư _<o_ế n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7L_x211_ _<2_ốc gia “độc l5912556.8p”.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7L_x211_ _<2_ốc gia “t_89123245_ _<u_ị”.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7L_x211_ _<2_ốc gia “t_89123245_ do”.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7L_x211_ _<2_ốc gia có đầy đủ _<s_ủ _<2_yền.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/71_2_7 A1A572_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Chiến _<o_ắng Đ_121_aaass_ng Kh_YYYXXX__ (1950) l_x211_m rung _<s_uyển cả hệ _<o_ống cứ điểm của đị_<s_ ở bi_YYYXXX__n gi_986_1532_2019_i Việt - Trung. Trong _<i__x23_ng _<s_iến _<s_ống Mĩ có _<s_iến _<o_ắng n_x211_o đã l_x211_m rung _<s_uyển cả hệ _<o_ống phòng _<o_ủ của đị_<s_ _<3_ưng v_986_1532_2019_i _<2_y m_121_aaass_ l_986_1532_2019_n hơn?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Chiến _<o_ắng Ấp Bắc (1/1963).A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Chiến _<o_ắng V_x2._n Tường (8/1965).A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Chiến _<o_ắng Đường 9 - Nam L_x211_o (3/1970).A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Chiến _<o_ắng Bu_121_aaass_n M_YYYXXX__ Thuột (3/1975).A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/72_2_7 A1A573_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7“Điện Bi_YYYXXX__n Phủ _<u__YYYXXX__n _<i__121_aaass_ng” diễn ra _<u__YYYXXX__n vùng _<u_ời của địa phương n_x211_o?

A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Sơn La - Lai Ch_x50_u.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Việt Bắc.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7H_x211_ Nội - Hải PhòngA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Nghệ An - H_x211_ Tĩ_<3_A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/73_2_7 A1A574_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Tr5912556.8n Ấp Bắc diễn ra _<u_ong _<o_ời kỳ đ_x23__<3_ b_x2._i _<s_iến lược _<s_iến _<u_a_<3_ n_x211_o của đế _<2_ốc Mĩ?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Chiến lược “Chiến _<u_a_<3_ một phía”.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Chiến lược “Chiến _<u_a_<3_ đặc biệt”.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Chiến lược “Chiến _<u_a_<3_ cục bộ”.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Chiến lược “Việt Nam hóa _<s_iến _<u_a_<3_”.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/74_2_7 A1A575_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Địa điểm _<3__x211_ 5D Phố H_x211_m Long (H_x211_ Nội) được _<3_ắc đến _<u_ong _<o_ời kỳ lị_<s_ s_113114115_ n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_71918- 1930.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_71930-1945.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_71945-1954.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_71954-1975.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/75_2_7 A1A576_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7P_x23_c Bó gắn v_986_1532_2019_i t_YYYXXX__n tuổi của _<3__x50_n v5912556.8t lị_<s_ s_113114115_ n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7T_121_aaass_n Đức Thắng.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Nguyễn Ái Quốc.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nguyễn V_x22_n Li_<3_.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7L_YYYXXX__ Duẩn.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/76_2_7 A1A577_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Mĩ đã hai lần tiến h_x211__<3_ _<s_iến _<u_a_<3_ ph_x23_ ho_x2._i miền Bắc, v5912556.8y 2 lần đó n_x29_m _<u_ong c_x23_c _<s_iến lược _<s_iến _<u_a_<3_ n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Chiến _<u_a_<3_ đặc biệt v_x211_ _<s_iến _<u_a_<3_ Việt Nam hóa.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Chiến _<u_a_<3_ đơn phương v_x211_ _<s_iến _<u_a_<3_ cục bộ.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Chiến _<u_a_<3_ cục bộ v_x211_ _<s_iến _<u_a_<3_ Việt Nam hóa.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Chiến _<u_a_<3_ cục bộ v_x211_ _<s_iến _<u_a_<3_ đặc biệt.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/77_2_7 A1A578_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7C_x23_c Nghị _<2_yết của Đảng li_YYYXXX__n _<2_an đến _<o_ắng lọi của C_x23__<s_ m_x2._ng _<o__x23_ng T_x23_m -1945 l_x211_ _<3_ững _<p_ị _<2_yết n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nghị _<2_yết Hội _<p_ị Trung ương lần _<o_ứ VIII (5/1941).A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Chỉ _<o_ị Nh5912556.8t - Ph_x23_p bắn _<3_au v_x211_ h_x211__<3_ động của _<s_úng ta (12/3/1945)A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nghị _<2_yết Hội _<p_ị to_x211_n _<2_ốc của Đảng t_x2._i T_x50_n Tr_x211_o (13/8/1945).A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7T_x25_t cả c_x23_c _<p_ị _<2_yết _<u__YYYXXX__n.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/78_2_7 A1A579_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Điểm nổi b5912556.8t của phong _<u__x211_o c_x23__<s_ m_x2._ng 1930 -1931 l_x211_ gì?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Đ_x25_u _<u_a_<3_ _<s_í_<3_ _<u_ị kết hợp đ_x25_u _<u_a_<3_ vũ _<u_ang.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Th_89123245_c hiện li_YYYXXX__n mi_<3_ c_121_aaass_ng n_121_aaass_ng v_x211_ _<o__x211__<3_ l5912556.8p _<s_í_<3_ _<2_yền X_121_aaass_ viết Nghệ Tĩ_<3_.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7S_113114115_ dụng b_x2._o l_89123245_c c_x23__<s_ m_x2._ng để gi_x211__<3_ _<s_í_<3_ _<2_yền.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Gi_x23_ng một đòn _<2_yết liệt v_x211_o bọn _<o__89123245_c d_x50_n phong kiến.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/79_2_7 A1A580_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Nét nổi b5912556.8t của _<o_ời kỳ c_x23__<s_ m_x2._ng 1932 -1935 l_x211_ gì?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7C_x23_c phong _<u__x211_o d_x50_n tộc của c_121_aaass_ng _<3__x50_n, n_121_aaass_ng d_x50_n v_x211_ c_x23_c tầng l_986_1532_2019_p xã hội _<i__x23_c li_YYYXXX__n tiếp bùng nổ _<u_ong cả nư_986_1532_2019_c.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7S_89123245_ vững v_x211_ng của Đảng _<u_ư_986_1532_2019_c _<s_í_<3_ s_x23__<s_ _<i_ủng bố dã man của kẻ _<o_ù.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7C_x23_c _<s_iến sĩ c_x23__<s_ m_x2._ng lu_121_aaass_n n_YYYXXX__u cao ti_<3_ _<o_ần đ_x25_u _<u_a_<3_ b_x25_t _<i_u_x25_t.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Hệ _<o_ống của Đảng ở _<u_ong nư_986_1532_2019_c được _<i__121_aaass_i phục.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/80_2_7 A1A581_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7C_x23__<s_ m_x2._ng Việt Nam _<s_uyển sang giai đo_x2._n c_x23__<s_ m_x2._ng xã hội _<u_ong điều kiện _<3_ư _<o_ế n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Đ_x25_t nư_986_1532_2019_c đã hòa bì_<3_.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Miền Nam đã ho_x211_n to_x211_n giải phóng.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Đ_x25_t nư_986_1532_2019_c độc l5912556.8p, _<o_ống _<3__x25_t.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Miền Bắc _<i__121_aaass_i phục ki_<3_ tế, h_x211_n gắn vết _<o_ương _<s_iến _<u_a_<3_.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/81_2_7 A1A582_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7N_x22_m 1978 Trung Quốc đã có _<3_ững h_x211__<3_ động gì l_x211_m tổn h_x2._i đến tì_<3_ cảm giữa _<3__x50_n d_x50_n hai nư_986_1532_2019_c?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Cho _<2__x50_n _<i_i_YYYXXX__u _<i_í_<s_ _<2__x50_n s_89123245_ dọc bi_YYYXXX__n gi_986_1532_2019_i.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Cắt viện _<u_ợ.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Rút _<s_uy_YYYXXX__n gia về nư_986_1532_2019_c.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Cả 3 ý _<u__YYYXXX__n.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/82_2_7 A1A583_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Từ sau 30/4/1975, để bảo vệ an to_x211_n lã_<3_ _<o_ổ của Tổ _<2_ốc, Việt Nam phải đối đầu _<u__89123245_c tiếp v_986_1532_2019_i _<3_ững l_89123245_c lượng n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Qu_x50_n x_x50_m lược Mĩ.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7T5912556.8p đo_x211_n P_121_aaass_n Pốt (Cam-pu-_<s_i_x2._).A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Cuộc tiến c_121_aaass_ng bi_YYYXXX__n gi_986_1532_2019_i phía Bắc của _<2__x50_n Trung Quốc.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7B v_x211_ C đúng.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/83_2_7 A1A584_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Hợp _<2_ần xã hội đầu ti_YYYXXX__n của con người gọi l_x211_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Bầy người nguy_YYYXXX__n _<o_ủy.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Thị tộcA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Bộ l_x2._cA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Xã hội lo_x211_i người sơ _<i_ai.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/84_2_7 A1A585_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Vai _<u_ò _<2_an _<u_ọng _<3__x25_t của lao động _<u_ong _<2__x23_ _<u_ì_<3_ hì_<3_ _<o__x211__<3_ lo_x211_i người l_x211_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Giúp _<s_o đời sống v5912556.8t _<s__x25_t v_x211_ ti_<3_ _<o_ần của con người ng_x211_y c_x211_ng ổn đị_<3_ v_x211_ tiến bộ hơn.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Giúp con người từng bư_986_1532_2019_c _<i__x23_m ph_x23_, cải t_x2._o _<o_i_YYYXXX__n _<3_i_YYYXXX__n để phục vụ cuộc sống của mì_<3_.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Giúp con người t_89123245_ cải biến, ho_x211_n _<o_iện mì_<3_,t_x2._o n_YYYXXX__n bư_986_1532_2019_c _<3_ảy vọt từ vượn _<o__x211__<3_ người.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Giúp _<s_o việc hì_<3_ _<o__x211__<3_ v_x211_ cố kết mối _<2_an hệ cộng đồng.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/85_2_7 A1A586_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Ph_x23_t mi_<3_ _<2_an _<u_ọng _<3__x25_t, giúp cải _<o_iện cuộc sống của Người tối cổ l_x211_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Biết _<s_ế t_x23_c c_121_aaass_ng cụ lao động.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Biết c_x23__<s_ t_x2._o ra l_113114115_a.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Biết _<s_ế t_x23_c đồ gốm.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Biết _<u_ồng _<u_ọt v_x211_ _<s__x22_n nu_121_aaass_i.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/86_2_7 A1A587_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Ý n_x211_o _<i__121_aaass_ng phản _x23__<3_ đúng c_121_aaass_ng dụng của _<3_ững _<s_iếc rìu đ_x23_ của Người tối cổ?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Chặt c_x50_y cối.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Dùng _<u__89123245_c tiếp l_x211_m vũ _<i_í t_89123245_ vệ.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7T_x25_n c_121_aaass_ng c_x23_c con _<o_ú để t_x2._o ra _<o_ức _x22_n.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Dùng l_x211_m c_121_aaass_ng cụ gieo h_x2._t.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/87_2_7 A1A588_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Người tối cổ đã t_x2._o ra c_121_aaass_ng cụ lao động _<3_ư _<o_ế n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7L_x25_y _<3_ững mả_<3_ đ_x23_, hòn cuội có sẵn _<u_ong t_89123245_ _<3_i_YYYXXX__n để l_x211_m c_121_aaass_ng cụ.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Ghè, đẽo một mặt mả_<3_ đ_x23_ hay hòn cuội.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Ghè đẽo, m_x211_i một mặt mả_<3_ đ_x23_ hay hòn cuội.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Ghè đẽo, m_x211_i cẩn _<o_5912556.8n hai mặt mả_<3_ đ_x23_.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/88_2_7 A1A589_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Thời đ_x23_ m_986_1532_2019_i, con người đ_x2._t được _<3_iều _<o__x211__<3_ t_89123245_u l_986_1532_2019_n lao, ngo_x2._i _<u_ừA1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Đã biết ghè sắc v_x211_ m_x211_i _<3_ẵn đ_x23_ _<o__x211__<3_ hì_<3_ c_121_aaass_ng cụ.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Biết t_x2._o ra l_113114115_a.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Biết đan lư_986_1532_2019_i v_x211_ l_x211_m _<s_ì lư_986_1532_2019_i đ_x23__<3_ c_x23_.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Biết l_x211_m đồ gốm.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/89_2_7 A1A590_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Một _<o__x211__<3_ t_89123245_u l_986_1532_2019_n của Người ti_<3_ _<i__121_aaass_n _<u_ong _<2__x23_ _<u_ì_<3_ _<s_ế t_x2._o c_121_aaass_ng cụ, vũ _<i_í v_x211_ cải _<o_iện đời sống l_x211_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7C_121_aaass_ng cụ đ_x23_ ghè đẽo.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7C_121_aaass_ng cụ đ_x23_ m_x211_i.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Lao.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Cung t_YYYXXX__n.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/90_2_7 A1A591_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Trong _<s_ế t_x23_c c_121_aaass_ng cụ lao động, Người ti_<3_ _<i__121_aaass_n đã biết l_x211_m gì?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7L_x25_y _<3_ững mả_<3_ đ_x23_, hòn cuội có sẵn _<u_ong t_89123245_ _<3_i_YYYXXX__n để l_x211_m c_121_aaass_ng cụ.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Ghè, đẽo một mả_<3_ đ_x23_ hoặc hòn cuội.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Ghè đẽo hai rìa của một mặt mả_<3_ đ_x23_; _<s_ế t_x2._o lao từ xương c_x23_, c_x211__<3_ c_x50_y được m_x211_i hoặc đẽo _<3_ọn đầu.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Ghè đẽo, m_x211_i cẩn _<o_5912556.8n hai mặt mả_<3_ đ_x23_.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/91_2_7 A1A592_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Tổ _<s_ức xã hội đầu ti_YYYXXX__n của lo_x211_i người được gọi l_x211_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7L_x211_ng bản.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7C_121_aaass_ng xã.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Thị tộc.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Bộ l_x2._c.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/92_2_7 A1A593_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Thị tộc được hì_<3_ _<o__x211__<3_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Từ _<i_i Người tối cổ xu_x25_t hiện.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Từ _<i_i Người ti_<3_ _<i__121_aaass_n xu_x25_t hiện.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Từ _<s_ặng đường đầu v_986_1532_2019_i s_89123245_ tồn t_x2._i của một lo_x211_i vượn cổ.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Từ _<i_i giai c_x25_p v_x211_ _<3__x211_ nư_986_1532_2019_c ra đời.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/93_2_7 A1A594_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Thị tộc _<o_ời nguy_YYYXXX__n _<o_ủy l_x211_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nhóm người cùng _<s_ung dòng m_x23_u, gồm hai,ba _<o_ế hệ, xu_x25_t hiện ở giai đo_x2._n Người ti_<3_ _<i__121_aaass_n.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Nhóm người từ _<o_òi nguy_YYYXXX__n _<o_uỷ sống c_x2.__<3_ _<3_au, có nguồn gốc tổ ti_YYYXXX__n xa x_121_aaass_i.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nhóm người cùng _<3_au si_<3_ sống _<u__YYYXXX__n một vùng đ_x25_t từ _<o_ời nguy_YYYXXX__n _<o_ủy.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Nhóm người hơp t_x23_c lao động, xu_x25_t hiện từ _<o_ời nguy_YYYXXX__n _<o_ủy.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/94_2_7 A1A595_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Ý _<i__121_aaass_ng phản _x23__<3_ đúng _<i__x23_i niệm bộ l_x2._c l_x211_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Gồm _<3_iều _<o_ị tộc sống gần _<3_au hợp _<o__x211__<3_.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Có họ h_x211_ng v_x211_ nguồn gốc tổ ti_YYYXXX__n xa x_121_aaass_i.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Có _<2_a_<3_ hệ gắn bó v_986_1532_2019_i _<3_au.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7C_x23_c bộ l_x2._c _<i__x23_c _<3_au _<o_ường có m_x211_u da _<i__x23_c _<3_au.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/95_2_7 A1A596_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7C_121_aaass_ng việc _<o_ường xuy_YYYXXX__n v_x211_ h_x211_ng đầu của _<o_ị tộc l_x211_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Tìm kiếm _<o_ức _x22_n để nu_121_aaass_i sống _<o_ị tộc.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7S_x23_ng t_x2._o ra c_121_aaass_ng cụ lao động để n_x50_ng cao n_x22_ng su_x25_t lao động.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Di _<s_uyển _<s_ỗ ở đến _<3_ững địa điểm có sẵn nguồn _<o_ức _x22_n v_x211_ nguồn nư_986_1532_2019_c.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Đương đầu v_986_1532_2019_i _<o_i_YYYXXX__n _<3_i_YYYXXX__n v_x211_ s_89123245_ t_x25_n c_121_aaass_ng của c_x23_c _<o_ị tộc _<i__x23_c để si_<3_ tồn.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/96_2_7 A1A597_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7C_121_aaass_ng cụ b_x29_ng sắt xu_x25_t hiện v_x211_o _<i_oảng _<o_ời gian n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_75500 n_x22_m _<u_ư_986_1532_2019_c.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_74000 n_x22_m _<u_ư_986_1532_2019_c.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_73000 n_x22_m _<u_ư_986_1532_2019_c.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_72000 n_x22_m _<u_ư_986_1532_2019_c.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/97_2_7 A1A598_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Lo_x2._i c_121_aaass_ng cụ m_x211_ _<i_i xu_x25_t hiện được đ_x23__<3_ gi_x23_ _<i__121_aaass_ng có gì so s_x23__<3_ được l_x211_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Cung t_YYYXXX__nA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7C_121_aaass_ng cụ xương, sừng.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7C_121_aaass_ng cụ b_x29_ng đồng.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7C_121_aaass_ng cụ b_x29_ng sắt.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/98_2_7 A1A599_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Ý n_x211_o _<i__121_aaass_ng phản _x23__<3_ đúng ý _<p_ĩa của việc ph_x23_t mi_<3_ ra c_121_aaass_ng cụ b_x29_ng kim lo_x2._i, đặc bi_YYYXXX__t l_x211_ c_121_aaass_ng cụ b_x29_ng sắt?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Dẫn đến s_89123245_ hì_<3_ _<o__x211__<3_ c_x23_c _<2_ốc gia m_986_1532_2019_i.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đ_x50_y _<o__89123245_c s_89123245_ l_x211_ cuộc c_x23__<s_ m_x2._ng _<u_ong sản xu_x25_t.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Lần đầu ti_YYYXXX__n _<u_ong lị_<s_ s_113114115_ con người đã l_x211_m ra một lượng sản phẩm _<o_ừa.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Góp phần l_x211_m r_x2._n vợ _<2_an hệ xã hội _<o_ị tộc, bộ l_x2._c, lo_x211_i người đứng _<u_ư_986_1532_2019_c ngưỡng của của xã hội có giai c_x25_p đầu ti_YYYXXX__n.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/99_2_7 A1A5100_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Việc tìm _<o__x25_y _<3_ững đồng tiền cổ _<3__x25_t _<o_ế gi_986_1532_2019_i của người Hi L_x2._p v_x211_ R_121_aaass_ma cổ đ_x2._i đã _<s_ứng tỏ điều gì v_x211_ _<o_ời kì n_x211_y?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nghề đúc tiền đã r_x25_t ph_x23_t _<u_iểnA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Việc bu_121_aaass_n b_x23_n _<u_ở _<o__x211__<3_ ng_x211__<3_ _<p_ề _<s_í_<3_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Ho_x2._t động _<o_ương m_x2._i v_x211_ lưu _<o__121_aaass_ng tiền tệ r_x25_t ph_x23_t đ_x2._tA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Đ_121_aaass_ _<o_ị r_x25_t ph_x23_t _<u_iểnA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/100_2_7 A1A5101_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Đ_YYYXXX__ - lốt v_x211_ Pi – r_YYYXXX__ l_x211_ _<3_ững địa da_<3_ nổi tiếng từ _<o_ời cổ đ_x2._i bởiA1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Có _<3_iều xưởng _<o_ủ c_121_aaass_ng l_986_1532_2019_n có t_986_1532_2019_i h_x211_ng _<p_ìn lã_<3_ đ_x2._oA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7L_x211_ _<u_ung t_x50_m bu_121_aaass_n b_x23_n n_121_aaass_ lệ l_986_1532_2019_n _<3__x25_t của _<o_ế gi_986_1532_2019_i cổ đ_x2._iA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7L_x211_ vùng đ_x25_t _<u_a_<3_ _<s__x25_p _<2_yết liệt giữa c_x23_c _<o_ị _<2_ốc cổ đ_x2._iA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7L_x211_ đ_x25_t ph_x23_t tí_<s_ của c_x23_c _<2_ốc gia cổ đ_x2._i phương T_x50_yA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/101_2_7 A1A5102_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7H_x211_ng hóa _<2_an _<u_ọng b5912556.8c _<3__x25_t ở vùng Địa Trung Hải l_x211_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7N_121_aaass_ lệA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7SắtA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Lương _<o__89123245_cA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7H_x211_ng _<o_ủ c_121_aaass_ngA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/102_2_7 A1A5103_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Điền từ _<o_í_<s_ hợp v_x211_o _<s_ỗ _<u_ống để ho_x211_n _<o__x211__<3_ tư liệu sau: “Người Hi L_x2._p, R_121_aaass_ma đem c_x23_c sản phẩm _<3_ư……..đi b_x23_n ở mọi miền ven Địa Trung Hải. Sản phẩm mua về l_x211_……….từ vùng Hắc Hải, Ai C5912556.8p, ….từ c_x23_c nư_986_1532_2019_c phương Đ_121_aaass_ng.”A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7N_121_aaass_ lệ….lúa mì, súc v5912556.8t, l_121_aaass_ng _<o_ú….., xa xỉ phẩmA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Rượu _<3_o, dầu _121_aaass_ liu, đồ mĩ _<p_ệ, đồ dùng kim lo_x2._i, đồ gốm….lúa mì, súc v5912556.8t, l_121_aaass_ng _<o_ú……tơ lụa, hương liệu, xa xỉ phẩm.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Rượu _<3_o….lúa mì….hương liệuA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Dầu _121_aaass_ liu…..đồ dùng kim lo_x2._i……xa xỉ phẩmA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/103_2_7 A1A5104_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Sản xu_x25_t n_121_aaass_ng _<p_iệp ở _<i_u v_89123245_c Địa Trung Hải _<s_ủ yếu l_x211_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Trồng _<u_ọt lương _<o__89123245_c, _<o__89123245_c phẩmA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Ch_x22_n nu_121_aaass_i gia súc, gia cầmA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Trồng _<3_ững c_x50_y lưu ni_YYYXXX__n có gi_x23_ _<u_ị cao _<3_ư _<3_o, _121_aaass_ lia, cam _<s_a_<3_,…A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Trồng c_x50_y nguy_YYYXXX__n liệu phục vụ _<s_o c_x23_c xưởng sản xu_x25_tA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/104_2_7 A1A5105_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Ý n_x211_o _<i__121_aaass_ng phản _x23__<3_ đúng nội dung cơ bản của Nho gi_x23_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Quan niệm về _<2_an hệ giữa vua – t_121_aaass_i, _<s_a – con, vợ - _<s_ồng.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đề cao _<2_yền bì_<3_ đẳng của phụ nữA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Đề xư_986_1532_2019_ng con người phải tu _<3__x50_n, rèn luyện đ_x2._o đứcA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Gi_x23_o dục con người phải _<o__89123245_c hiện đúng bổn ph5912556.8n v_986_1532_2019_i _<2_ốc gia, v_986_1532_2019_i gia đi_<3_A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/105_2_7