A1A5_x2905__2_7x12515x185x125x1765x12055x11065x15x11535x1755x12415x11825x165x1315x1505x12525x11755A1A5/_x2905__2_7A1A5_..rt)(dfdf)_----_2_7A1A5_01rtfg_-_dg.__d-gdg_2_7Lị_<s_ S_113114115_ 6A1A5/_01rtfg_-_dg.__d-gdg_2_7A1A5ghi_<s_u_2_7Ôn T5912556.8p Lị_<s_ S_113114115_ 6 (Tổng hợp)A1A5/ghi_<s_u_2_7A1A5/_..rt)(dfdf)_----_2_7A1A5t_uD_R_2_7A1A5/t_uD_R_2_7
 A1A50_2_7A1A5_anti_vs_xem__2_7B_x29_ng kiến _<o_ức đã học em hãy _<s_o biết lị_<s_ s_113114115_ l_x211_ gì? A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Những gì đang diễn raA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Những gì _<s_ưa diễn raA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Những gì sẽ diễn raA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Những gì đã diễn ra _<u_ong _<2__x23_ _<i_ứA1A5/_0x001520_4_2_7A1A5/0_2_7 A1A51_2_7A1A5_anti_vs_xem__2_7Lị_<s_ s_113114115_ lo_x211_i người l_x211_?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Tìm hiểu _<3_ững ho_x2._t động của con người hiện nayA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7D_89123245_ng l_x2._i ho_x2._t động của con người, xã hội lo_x211_i người từ _<i_i xu_x25_t hiện đến nayA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Tìm hiểu ho_x2._t động của xã hội lo_x211_i người hiện nayA1A5/_0x001520_3_2_7A1A5/1_2_7 A1A52_2_7A1A5_anti_vs_xem__2_7Học lị_<s_ s_113114115_ để l_x211_m gì?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Biết _<s_o vuiA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7T_121_aaass_ điểm _<s_o cuộc sốngA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Hiểu cội nguồn của tổ ti_YYYXXX__n, _<s_a _121_aaass_ngA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Biết việc l_x211_m của người xưaA1A5/_0x001520_4_2_7A1A5/2_2_7 A1A53_2_7A1A5_anti_vs_xem__2_7C_x50_u da_<3_ ng_121_aaass_n "Lị_<s_ s_113114115_ l_x211_ _<o_ầy d_x2._y của cuộc sống" l_x211_ của ai?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7L_YYYXXX__ NinA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Xi X_YYYXXX__ R_121_aaass_ngA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7B_x23_c HồA1A5/_0x001520_3_2_7A1A5/3_2_7 A1A54_2_7A1A5_anti_vs_xem__2_7Để hiểu biết lị_<s_ s_113114115_, ta d_89123245_a v_x211_o:A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Tư liệu _<u_uyền miệng, hiện v5912556.8t, _<s_ữ viếtA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đồ v5912556.8tA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Bản đồA1A5/_0x001520_3_2_7A1A5/4_2_7 A1A55_2_7A1A5_anti_vs_xem__2_7Tư liệu hiện v5912556.8t gồm:A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Di tí_<s_ đồ v5912556.8t của người xưaA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Lời kểA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7C_x50_u _<s_uyệnA1A5/_0x001520_3_2_7A1A5/5_2_7 A1A56_2_7A1A5_anti_vs_xem__2_7Tư liệu _<s_ữ biết gồmA1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Đồ v5912556.8tA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Hì_<3_ ả_<3_A1A5/_0x001520_2_2_7A1A5/6_2_7 A1A57_2_7A1A5_anti_vs_xem__2_7Di tí_<s_ lị_<s_ s_113114115_ của Phú Thọ l_x211_?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Th_x211__<3_ Cổ LoaA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đền hùngA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7V_x22_n Miếu Quốc T_113114115_ Gi_x23_m.A1A5/_0x001520_3_2_7A1A5/7_2_7 A1A58_2_7A1A5_anti_vs_xem__2_7C_x50_u da_<3_ ng_121_aaass_n "Lị_<s_ s_113114115_ l_x211_ _<o_ầy d_x2._y của cuộc sống" em hiểu c_x50_u _x25_y _<3_ư _<o_ế n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Cung c_x25_p b_x211_i học lị_<s_ s_113114115_ _<s_o người đời sauA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Người đời nay cần biết s_113114115_A1A5/_0x001520_2_2_7A1A5/8_2_7 A1A59_2_7A1A5_anti_vs_xem__2_7Lị_<s_ s_113114115_ cần x_x23_c đị_<3_ _<o_ời gian vì:A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Thời gian l_x211_ v_x211_ng ngọcA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7C_x23_c s_89123245_ kiện xảy ra ở _<o_ời gian _<3__x25_t đị_<3_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Muốn tìm hiểu v_x211_ d_89123245_ng l_x2._i lị_<s_ s_113114115_ _<o_ì cần phải sắp xếp c_x23_c s_89123245_ kiện đó _<o_eo _<o_ứ t_89123245_ _<o_ời gianA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7S_89123245_ kiện cần có tuổiA1A5/_0x001520_4_2_7A1A5/9_2_7 A1A510_2_7A1A5_anti_vs_xem__2_7Để tí_<3_ _<o_ời gian, con người đã d_89123245_a v_x211_i:A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Á_<3_ s_x23_ngA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Thời tiếtA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Mùa vụA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Chu kỳ mọc, lặn, di _<s_uyển của mặt _<u_ời, mặt _<u__x22_ng.A1A5/_0x001520_4_2_7A1A5/10_2_7 A1A511_2_7A1A5_anti_vs_xem__2_7Âm Lị_<s_ l_x211_?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Di _<s_uyển của _<u__x23_i đ_x25_tA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Di _<s_uyển của mặt _<u_ờiA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Di _<s_uyển của c_x23_c vì saoA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Tí_<3_ _<o_eo s_89123245_ di _<s_uyển mặt _<u__x22_ng _<2_a_<3_ _<u__x23_i đ_x25_tA1A5/_0x001520_4_2_7A1A5/11_2_7 A1A512_2_7A1A5_anti_vs_xem__2_7Dương lị_<s_ l_x211_?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Tí_<3_ _<o_eo di _<s_uyển của mặt _<u_ờiA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Di _<s_uyển của _<u__x23_i đ_x25_tA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Tí_<3_ _<o_eo s_89123245_ di _<s_uyển của _<u__x23_i đ_x25_t _<2_a_<3_ mặt _<u_ờiA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Di _<s_uyển sao hỏaA1A5/_0x001520_4_2_7A1A5/12_2_7 A1A513_2_7A1A5_anti_vs_xem__2_7Vì sao _<o_ế gi_986_1532_2019_i cần một _<o_ứ lị_<s_ _<s_ung:A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Nhu cầu một nư_986_1532_2019_cA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Nhu cầu con ngườiA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nhu cầu bu_121_aaass_n b_x23_nA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Nhu cầu giao lưu c_x23_c nư_986_1532_2019_c, c_x23_c _<i_u v_89123245_c cần _<o_ống _<3__x25_t c_x23__<s_ tí_<3_.A1A5/_0x001520_4_2_7A1A5/13_2_7 A1A514_2_7A1A5_anti_vs_xem__2_7C_121_aaass_ng lị_<s_ được tí_<3_:A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7L_x25_y n_x22_m tương _<u_uyền _<s_úa Gi_YYYXXX__ Xu ra đời l_x211_ n_x22_m đầu ti_YYYXXX__n của c_121_aaass_ng nguy_YYYXXX__n.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_x22_m ra đời của X_YYYXXX__ DaA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7N_x22_m ra đời của Pom P_YYYXXX__A1A5/_0x001520_3_2_7A1A5/14_2_7 A1A515_2_7A1A5_anti_vs_xem__2_7N_x22_m 179 TCN hiểu l_x211_:A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7C_x23__<s_ hiện nay l_x211_ 179 n_x22_mA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_72000 n_x22_mA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7C_x23__<s_ 179 n_x22_m m_986_1532_2019_i đến n_x22_m đầu CNA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_72179 n_x22_mA1A5/_0x001520_4_2_7A1A5/15_2_7 A1A516_2_7A1A5_anti_vs_xem__2_7Một _<o_i_YYYXXX__n ni_YYYXXX__n kỷ gồm bao _<3_i_YYYXXX__u n_x22_m?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_71000 n_x22_mA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7100 n_x22_mA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_710 n_x22_mA1A5/_0x001520_3_2_7A1A5/16_2_7 A1A517_2_7A1A5_anti_vs_xem__2_7N_x22_m 201 _<o_uộc _<o_ế kỷ m_x25_y?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Thế kỷ IIIA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Thế Kỷ IVA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Thế Kỉ IIA1A5/_0x001520_3_2_7A1A5/17_2_7 A1A518_2_7A1A5_anti_vs_xem__2_7C_x23__<s_ tí_<3_ _<i_oảng _<o_ời gian của s_89123245_ kiện: Nư_986_1532_2019_c Âu L_x2._c bị Tri_YYYXXX__u Đ_x211_ x_x50_m _<s_iếm 179 _<u_ư_986_1532_2019_c c_121_aaass_ng nguy_YYYXXX__n đến n_x22_m 2004?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_72004 - 179 = 1825A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_72002 n_x22_mA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_72004 + 179 = 2183 n_x22_mA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7179 n_x22_mA1A5/_0x001520_4_2_7A1A5/18_2_7 A1A519_2_7A1A5_anti_vs_xem__2_7Qu_YYYXXX__ hương của phong _<u__x211_o v_x22_n hóa Phục Hưng l_x211_ nư_986_1532_2019_c n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Nư_986_1532_2019_c Ph_x23_pA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Nư_986_1532_2019_c BỉA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nư_986_1532_2019_c A_<3_A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Nư_986_1532_2019_c ÝA1A5/_0x001520_4_2_7A1A5/19_2_7 A1A520_2_7A1A5_anti_vs_xem__2_7Giữa _<o_ế kỉ XIX, hầu hết c_x23_c _<2_ốc gia Đ_121_aaass_ng Nam Á đều _<u_ở _<o__x211__<3_ _<o_uộc địa của _<s_ủ _<p_ĩa _<o__89123245_c d_x50_n phương T_x50_y, _<u_ừ nư_986_1532_2019_c n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Việt NamA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Th_x23_i LanA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Phi-lip-pinA1A5/_0x001520_3_2_7A1A5/20_2_7 A1A521_2_7A1A5_anti_vs_xem__2_7L_89123245_c lượng sản xu_x25_t _<s_ủ yếu _<u_ong c_x23_c lã_<3_ địa phong kiến l_x211_ ai?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7N_121_aaass_ng d_x50_n t_89123245_ doA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_121_aaass_ng _<o__121_aaass_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7N_121_aaass_ lệA1A5/_0x001520_3_2_7A1A5/21_2_7 A1A522_2_7A1A5_anti_vs_xem__2_7Để dẹp “Lo_x2._n 12 sứ _<2__x50_n”, Đi_<3_ Bộ Lĩ_<3_ đã li_YYYXXX__n kết v_986_1532_2019_i:A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Sứ _<2__x50_n Trần LãmA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Sứ _<2__x50_n Nguyễn Thủ TiệpA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Sứ _<2__x50_n Ng_121_aaass_ Nh5912556.8t Kh_x23__<3_A1A5/_0x001520_3_2_7A1A5/22_2_7 A1A523_2_7A1A5_anti_vs_xem__2_7Đi_<3_ Bộ Lĩ_<3_ được _<3__x50_n d_x50_n t_121_aaass_n xưng l_x211_:A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Bắc Bì_<3_ VươngA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Bì_<3_ Đi_<3_ VươngA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Bố C_x23_i Đ_x2._i VươngA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7V_x2._n Thắng VươngA1A5/_0x001520_4_2_7A1A5/23_2_7 A1A524_2_7A1A5_anti_vs_xem__2_7Nguy_YYYXXX__n _<3__x50_n n_x211_o dư_986_1532_2019_i đ_x50_y đã giúp Đi_<3_ Bộ Lĩ_<3_ _<o_ống _<3__x25_t dược đ_x25_t nư_986_1532_2019_c?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7S_89123245_ ủng hộ của _<3__x50_n d_x50_nA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7T_x211_i n_x22_ng của Đị_<3_ Bộ Lĩ_<3_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7S_89123245_ li_YYYXXX__n kết của c_x23_c sứ _<2__x50_nA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7T_x25_t cả c_x23_c ý _<u__YYYXXX__nA1A5/_0x001520_4_2_7A1A5/24_2_7 A1A525_2_7A1A5_anti_vs_xem__2_7Trong ho_x211_n cả_<3_ lị_<s_ s_113114115_ n_x211_o L_YYYXXX__ Ho_x211_n l_YYYXXX__n ng_121_aaass_i Ho_x211_ng đế?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Nội bộ _<u_iều đì_<3_ m_x50_u _<o_uẫn sau _<i_i Đi_<3_ Ti_YYYXXX__n Ho_x211_n m_x25_tA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đi_<3_ Ti_YYYXXX__n Ho_x211_ng m_x25_t, vua kết vị còn _<3_ỏ, _<3__x211_ Tống _<s_uẩn bị x_x50_m lược nư_986_1532_2019_c ta.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Thế l_89123245_c L_YYYXXX__ Ho_x211_n m_x2.__<3_, ép _<3__x211_ Đi_<3_ _<3_ường ng_121_aaass_i.A1A5/_0x001520_3_2_7A1A5/25_2_7 A1A526_2_7A1A5_anti_vs_xem__2_7Dư_986_1532_2019_i _<o_ời _<3__x211_ Lý, đến n_x22_m 1054, Quốc hiệu nư_986_1532_2019_c ta l_x211_ gì?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Đ_x2._i ViệtA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đ_x2._i Cồ ViệtA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Đ_x2._i NamA1A5/_0x001520_3_2_7A1A5/26_2_7 A1A527_2_7A1A5_anti_vs_xem__2_7V_x211_o _<o_ời gian n_x211_o _<2__x50_n Tống vượt ải Nam Quan _<2_a L_x2._ng Sơn tiến v_x211_o nư_986_1532_2019_c ta?                                                                                               A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Cuối n_x22_m 1076A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Cuối n_x22_m 1075A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Đầu n_x22_m 1077A1A5/_0x001520_3_2_7A1A5/27_2_7 A1A528_2_7A1A5_anti_vs_xem__2_7Chùa Một Cột ở H_x211_ Nội được x_x50_y d_89123245_ng v_x211_o _<o_ời n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7Thời Tiền L_YYYXXX__A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Thời TrầnA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Thời H5912556.8u L_YYYXXX__A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Thời LýA1A5/_0x001520_4_2_7A1A5/28_2_7 A1A529_2_7A1A5_anti_vs_xem__2_7V_x22_n Miếu được x_x50_y d_89123245_ng v_x211_o n_x22_m n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5_0x001520_1_2_7N_x22_m 1075A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_x22_m 1070A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7N_x22_m 1080A1A5/_0x001520_3_2_7A1A5/29_2_7 A1A530_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Nh_x211_ Trần huy động _<3__x50_n d_x50_n cả nư_986_1532_2019_c đắp đ_YYYXXX__ dọc hai bờ c_x23_c con s_121_aaass_ng l_986_1532_2019_n v_x211_o n_x22_m n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7N_x22_m 1225A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_x22_m 1252A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7N_x22_m 1247A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7N_x22_m 1248A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/30_2_7 A1A531_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7T_x23_c phẩm “Bi_<3_ _<o_ư yếu lược” do ai viết?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Trần Quang KhảiA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Trần Quốc Tu_x25_nA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Trần Hưng Đ_x2._oA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Trần Nguy_YYYXXX__n Đ_x23_nA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/31_2_7 A1A532_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Người n_x211_o đã d_x50_ng s_986_1532_2019_ đòi vua _<s_ém đầu 7 t_YYYXXX__n nị_<3_ _<o_ần?   A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nguyễn Phi Kha_<3_A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Trần Quốc Tu_x25_nA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Trần Kh_x23__<3_ DưA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Chu V_x22_n AnA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/32_2_7 A1A533_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Giai c_x25_p tư sản _<s__x50_u Âu được hì_<3_ _<o__x211__<3_ từ tầng l_986_1532_2019_p n_x211_o dư_986_1532_2019_i đ_x50_y?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Địa _<s_ủ gi_x211_u cóA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Thương _<3__x50_n gi_x211_u cóA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Chủ xưởng, _<s_ủ đồn điềnA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7C_x50_u B v_x211_ C đúngA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/33_2_7 A1A534_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Điền từ còn _<o_iếu v_x211_o _<s_ỗ _<u_ống _<u_ong c_x50_u sau:
... góp phần _<o_úc đẩy _<o_ương _<p_iệp _<s__x50_u Âu ph_x23_t _<u_iển v_x211_ đem l_x2._i _<s_o giai c_x25_p tư sản _<s__x50_u Âu _<3_ững nguồn nguy_YYYXXX__n liệu _<2_ý gi_x23_, _<3_ững vùng đ_x25_t m_YYYXXX___<3_ m_121_aaass_ng ở _<s__x50_u Á, _<s__x50_u Phi v_x211_ _<s__x50_u Mĩ.
A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7S_89123245_ xu_x25_t hiện của _<o__x211__<3_ mịA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Cuộc ph_x23_t kiến địa líA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Những _<s_uyến đi biển vòng _<2_a_<3_ _<o_ế gi_986_1532_2019_iA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7T_x25_t cả đều đúngA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/34_2_7 A1A535_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Giai c_x25_p tư sản đang l_YYYXXX__n ở _<s__x50_u Âu đã _<s_ống l_x2._i hệ tư tưởng của t_121_aaass_n gi_x23_o n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Hồi gi_x23_oA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Ki-t_121_aaass_ gi_x23_oA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Ph5912556.8t gi_x23_oA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Ấn độ gi_x23_oA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/35_2_7 A1A536_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7 “Lo_x2._n 12 sứ _<2__x50_n” diễn ra _<u_ong _<o_ời điểm lị_<s_ s_113114115_ n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Cuối _<o_ời Đi_<3_A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đầu _<o_ời Đi_<3_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Cuối _<o_ời Ng_121_aaass_A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Đầu _<o_ời Ng_121_aaass_A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/36_2_7 A1A537_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Cơ c_x25_u h_x211__<3_ _<s_í_<3_ dư_986_1532_2019_i _<o_ời _<3__x211_ Lý được sắp xếp _<o_eo _<o_ứ t_89123245_ n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Lộ - Huyện - Hương, xãA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Lộ - Phủ - Ch_x50_u - Hương, xãA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Lộ - Phủ - Ch_x50_u, xãA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Lộ - Phủ - Huyện - Hương, xãA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/37_2_7 A1A538_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Nguy_YYYXXX__n tắc m_x211_ _<3__x211_ Lý lu_121_aaass_n ki_YYYXXX__n _<2_yết giữ vững _<u_ong _<i_i duy _<u_ì mối giao bang v_986_1532_2019_i c_x23_c nư_986_1532_2019_c l_x23_ng giềng l_x211_:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Hòa hảo, _<o__x50_n _<o_iệnA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đo_x211_n kết, _<u__x23__<3_ xung độtA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Mở c_113114115_a, _<u_ao đổi, lưu _<o__121_aaass_ng h_x211_ng hóaA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Giữ vững _<s_ủ _<2_yền v_x211_ to_x211_n vẹn lã_<3_ _<o_ổA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/38_2_7 A1A539_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Tì_<3_ hì_<3_ ki_<3_ tế, xã hội Việt Nam _<3_ững n_x22_m 60 của _<o_ế kỉ XIX _<3_ư _<o_ế n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Ki_<3_ tế, xã hội _<i_ủng hoảng _<p_i_YYYXXX__m _<u_ọng.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_121_aaass_ng _<p_iệp, _<o_ủ c_121_aaass_ng _<p_iệp, _<o_ương _<p_iệp đì_<3_ _<u_ệ.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7M_x50_u _<o_uẫn giai c_x25_p v_x211_ m_x50_u _<o_uẫn d_x50_n tộc gay gắt.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7T_x211_i _<s_í_<3_ c_x2._n kiệt, _<3__x50_n d_x50_n đói _<i_ổ.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/39_2_7 A1A540_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Cuộc _<i_ởi _<p_ĩa của bi_<3_ lí_<3_ v_x211_ d_x50_n phu n_x22_m 1866 dư_986_1532_2019_i s_89123245_ _<o_am gia của một số sĩ phu, _<2_an l_x2._i _<2_ý tộc nổ ra ở đ_x50_u?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Huế                    A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Bắc Ni_<3_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Tuy_YYYXXX__n QuangA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Th_x23_i Nguy_YYYXXX__nA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/40_2_7 A1A541_2_7A1A5_anti_vs_xem__2_7S_x23__<s_ Lị_<s_ s_113114115_ 8 _<u_ang 134: N_YYYXXX__u _<3_ững _<3_5912556.8n xét _<s_í_<3_ về tì_<3_ hì_<3_ ki_<3_ tế, xã hội Việt Nam giữa _<o_ế kỉ XIX.A1A5/_anti_vs_xem__2_7A1A5_pass_15x_091__2_7Giữa _<o_ế kỉ XIX, nền ki_<3_ tế-xã hội Việt Nam rơi v_x211_o tì_<3_ _<u__x2._ng _<i_ủng hoảng _<p_i_YYYXXX__m _<u_ọng: Bộ m_x23_y _<s_í_<3_ _<2_yền từ _<u_ung ương đến địa phương mục ruỗng, n_121_aaass_ng _<p_iệp, _<o_ủ c_121_aaass_ng _<p_iệp v_x211_ _<o_ương _<p_iệp sa sút, t_x211_i _<s_í_<3_ _<i__121_aaass_ kiệt, đời sống _<3__x50_n d_x50_n v_121_aaass_ cùng _<i_ó _<i__x22_n, m_x50_u _<o_uẫn giai c_x25_p v_x211_ m_x50_u _<o_uẫn xã hội ng_x211_y c_x211_ng gay gắt l_x211_m _<s_o xã hội _<o__YYYXXX__m rối lo_x2._n.A1A5/_pass_15x_091__2_7A1A5/41_2_7 A1A542_2_7 A1A5_anti_vs_xem__2_7Lị_<s_ s_113114115_ l_986_1532_2019_p 8 _<u_ang 134 SGK: Nguy_YYYXXX__n _<3__x50_n n_x211_o dẫn đến _<3_ững cuộc _<i_ởi _<p_ĩa n_121_aaass_ng d_x50_n _<s_ống _<u_iều đì_<3_ phong kiến _<u_ong n_113114115_a cuối _<o_ế kỉ XIX?A1A5/_anti_vs_xem__2_7 A1A5_pass_15x_091__2_7Bộ m_x23_y _<s_í_<3_ _<2_yền mục m_x23_t từ _<u_ung ương đến địa phương, ki_<3_ tế sa sút, _<3__x50_n d_x50_n bị _x23_p bức một cổ hai _<u_òng (s_89123245_ bóc lột của _<u_iều đì_<3_ phong kiến, s_89123245_ bóc lột đ_x211_n _x23_p của _<s_í_<3_ _<2_yền đ_121_aaass_ hộ), đời sống v_121_aaass_ cùng c_89123245_c _<i_ổ =_2_7 phong _<u__x211_o _<i_ởi _<p_ĩa của n_121_aaass_ng d_x50_n l_x2._i tiếp tục bùng nổ dữ dội _<u_ong _<3_ững n_x22_m cuối _<o_ế kỉ XIX.A1A5/_pass_15x_091__2_7A1A5/42_2_7 A1A543_2_7 A1A5_anti_vs_xem__2_7Lị_<s_ s_113114115_ l_986_1532_2019_p 8 _<u_ang 135 SGK: Vì sao c_x23_c _<2_an l_x2._i, sĩ phu đưa ra _<3_ững đề _<p_ị cải c_x23__<s_?A1A5/_anti_vs_xem__2_7 A1A5_pass_15x_091__2_7- Đ_x25_t nư_986_1532_2019_c đang _<u_ong tì_<3_ _<u__x2._ng nguy _<i_ốn (Ph_x23_p mở rộng x_x50_m lược; _<u_iều đì_<3_ bảo _<o_ủ, l_x2._c h5912556.8u: Ki_<3_ tế kiệt _<2_ệ; m_x50_u _<o_uẫn xã hội gay gắt...).

- Xu_x25_t ph_x23_t từ lòng y_YYYXXX__u nư_986_1532_2019_c.

- C_x23_c sĩ phu l_x211_ _<3_ững người _<o__121_aaass_ng _<o__x23_i, đi _<3_iều, biết _<3_iều, đã từng được _<s_ứng kiến s_89123245_ phồn _<o_ị_<3_ của tư bản Âu - Mĩ v_x211_ _<o__x211__<3_ t_89123245_u của nền v_x22_n ho_x23_ phương T_x50_y.A1A5/_pass_15x_091__2_7A1A5/43_2_7 A1A544_2_7 A1A5_anti_vs_xem__2_7Lị_<s_ s_113114115_ l_986_1532_2019_p 8 _<u_ang 135 SGK: Kể t_YYYXXX__n _<3_ững sĩ phu ti_YYYXXX__u biểu _<u_ong phong _<u__x211_o cải c_x23__<s_ ở n_113114115_a cuối _<o_ế kỉ XIX. N_YYYXXX__u _<3_ững nội dung _<s_í_<3_ _<u_ong c_x23_c đề _<p_ị cải c_x23__<s_ của họ.A1A5/_anti_vs_xem__2_7 A1A5_pass_15x_091__2_7- Trần Đì_<3_ Túc v_x211_ Nguyễn Huy Tế (1868): Xin mở c_113114115_a biển Tr_x211_ Lí (Nam Đị_<3_).

- Đi_<3_ V_x22_n Điền (1868) xin đẩy m_x2.__<3_ việc _<i_ai _<i_ẩn đ_x25_t hoang v_x211_ _<i_ai mỏ, ph_x23_t _<u_iển bu_121_aaass_n b_x23_n, _<s__x25_n _<s_ỉ_<3_ _<2_ốc phòng.

- Nguyễn Trường Tộ (1863 - 1871): Đề _<p_ị _<s__x25_n _<s_ỉ_<3_ bộ m_x23_y _<2_an l_x2._i, ph_x23_t _<u_iển c_121_aaass_ng, _<o_ương _<p_iệp v_x211_ t_x211_i _<s_í_<3_, _<s_ỉ_<3_ đốn võ bị, mở rộng ngo_x2._i giao, cải tổ gi_x23_o dục.

- Nguyễn Lộ Tr_x2.__<s_ (1877-1882): Đề _<p_ị _<s__x25_n hưng d_x50_n _<i_í, _<i_ai _<o__121_aaass_ng d_x50_n _<u_í, bảo vệ đ_x25_t nư_986_1532_2019_c.A1A5/_pass_15x_091__2_7A1A5/44_2_7 A1A545_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7 Đầu _<o_ế kỉ XX, đứng đầu Nh_x211_ nư_986_1532_2019_c _<2__x211_n _<s_ủ _<s_uy_YYYXXX__n _<s_ế ở Nga l_x211_ ai?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nga ho_x211_ng Ni-c_121_aaass_-lai I.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Nga ho_x211_ng Ni-c_121_aaass_-lai II.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nga ho_x211_ng Ni-c_121_aaass_-lai III.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Nga Ho_x211_ng Đ_x2._i ĐếA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/45_2_7 A1A546_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Nga ho_x211_ng _<o_am gia Chiến _<u_a_<3_ _<o_ế gi_986_1532_2019_i _<o_ứ _<3__x25_t (1914 - 1918) đã đẩy nư_986_1532_2019_c Nga v_x211_o tì_<3_ _<u__x2._ng:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Khủng hoảng _<u_ầm _<u_ọng về ki_<3_ tế.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_x2._n _<o__x25_t _<p_iệp t_x22_ng _<3_a_<3_, n_x2._n đói xảy ra _<u_ầm _<u_ọngA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Khủng hoảng _<u_ầm _<u_ọng về ki_<3_ tế, _<s_í_<3_ _<u_ị - xã hội.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Bị c_x23_c nư_986_1532_2019_c đế _<2_ốc _<o__121_aaass_n tí_<3_.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/46_2_7 A1A547_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Tì_<3_ hì_<3_ nư_986_1532_2019_c Nga _<u_ư_986_1532_2019_c _<i_i c_x23__<s_ m_x2._ng bùng nổ?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7L_x211_ một đế _<2_ốc _<2__x50_n _<s_ủ _<s_uy_YYYXXX__n _<s_ế bảo _<o_ủ về _<s_í_<3_ _<u_ị, l_x2._c h5912556.8u về ki_<3_ tế.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7H5912556.8u _<2_ả của cuộc _<s_iến _<u_a_<3_ (1914) đè nặng l_YYYXXX__n c_x23_c tầng l_986_1532_2019_p _<3__x50_n d_x50_n đặc biệt l_x211_ n_121_aaass_ng d_x50_n, m_x50_u _<o_uẫn xã hội ph_x23_t _<u_iển gay gắt.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Chí_<3_ phủ Nga ho_x211_ng b_x25_t l_89123245_c, _<i__121_aaass_ng còn _<i_ả n_x22_ng tiếp tục _<o_ống _<u_ị.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7T_x25_t cả c_x23_c ý _<u__YYYXXX__n.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/47_2_7 A1A548_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7H5912556.8u _<2_ả _<p_i_YYYXXX__m _<u_ọng _<3__x25_t nư_986_1532_2019_c Nga g_x23__<3_ _<s_ịu do _<s_i_YYYXXX__n _<u_a_<3_ đế _<2_ốc (1914-1918) để l_x2._i :A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Ki_<3_ tế suy sụp.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Li_YYYXXX__n tiếp _<o_ua _<u_5912556.8n, xã hội _<i__121_aaass_ng ổn đị_<3_.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Ki_<3_ tế suy sụp, _<2__x50_n đội _<o_iếu vũ _<i_í lương _<o__89123245_c.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Ki_<3_ tế suy sụp, m_x50_u _<o_uẫn xã hội gay gắt.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/48_2_7 A1A549_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Vì sao _<3__x50_n d_x50_n _<s__x23_n ghét Nga ho_x211_ng ?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nga ho_x211_ng bóc lột _<3__x50_n d_x50_n _<o__x50_m tệ.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Nga ho_x211_ng đẩy _<3__x50_n d_x50_n Nga v_x211_o cuộc _<s_iến _<u_a_<3_ đế _<2_ốcA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nga ho_x211_ng đ_x23__<3_ _<o_uế ruộng đ_x25_t cao.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Nga ho_x211_ng _<i__121_aaass_ng _<u_ang bị đầy đủ vũ _<i_í _<s_o _<2__x50_n đội.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/49_2_7 A1A550_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Đầu _<o_ế kỉ XX, nư_986_1532_2019_c Nga đứng _<u_ư_986_1532_2019_c một tì_<3_ _<o_ế _<3_ư _<o_ế n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Bùng nổ cuộc c_x23__<s_ m_x2._ng để xóa bỏ _<s_ế độ Nga ho_x211_ng.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7C_x23_c nư_986_1532_2019_c đế _<2_ốc lần lượt _<o__121_aaass_n tí_<3_ Nga.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Chí_<3_ phủ Nga ho_x211_ng sắp bị sụp đổ.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Ki_<3_ tế bị _<i_ủng hoảng _<u_ầm _<u_ọng.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/50_2_7 A1A551_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Phải l5912556.8t đổ _<s_í_<3_ phủ Nga ho_x211_ng để tổ _<s_ức nư_986_1532_2019_c Cộng hòa d_x50_n _<s_ủ Nga, _<o__89123245_c hiện ng_x211_y l_x211_m 8 giờ v_x211_ _<u_ao to_x211_n bộ ruộng đ_x25_t _<s_o n_121_aaass_ng d_x50_n. Đó l_x211_ lời k_YYYXXX__u gọi của tổ _<s_ức n_x211_o ?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Ban _<s__x25_p h_x211__<3_ Đảng bộ P_YYYXXX__-tơ-r_121_aaass_-gr_x23_t.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đảng C_121_aaass_ng _<3__x50_n Xã hội d_x50_n _<s_ủ Nga.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Quốc tế _<o_ứ _<3__x25_t.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Quốc tế _<o_ứ hai.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/51_2_7 A1A552_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7L_89123245_c lượng _<o_am gia C_x23__<s_ m_x2._ng _<o__x23_ng Hai-1917 ở Nga l_x211_ :A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Phụ nữ, n_121_aaass_ng d_x50_n.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Phụ nữ, c_121_aaass_ng _<3__x50_n, bi_<3_ lí_<3_A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Phụ nữ, c_121_aaass_ng _<3__x50_n, n_121_aaass_ng d_x50_n.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7 C_121_aaass_ng _<3__x50_n, n_121_aaass_ng d_x50_n.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/52_2_7 A1A553_2_7 A1A5_anti_vs_xem__2_7Vì sao sau _<i_i C_x23__<s_ m_x2._ng _<o__x23_ng Hai _<o__x211__<3_ c_121_aaass_ng, L_YYYXXX__-nin v_x211_ Đảng B_121_aaass_n-s_YYYXXX__-ví_<s_ phải _<s_uẩn bị kế ho_x2.__<s_ tiếp tục l_x211_m c_x23__<s_ m_x2._ng? A1A5/_anti_vs_xem__2_7 A1A5_pass_15x_091__2_7- C_x23__<s_ m_x2._ng d_x50_n _<s_ủ tư sản _<o__x23_ng Hai 1917 tuy đã l5912556.8t đổ _<s_ế độ Nga ho_x211_ng, _<o__89123245_c hiện _<o__x211__<3_ c_121_aaass_ng một phần của _<3_iệm vụ c_x23__<s_ m_x2._ng tư sản, song ở nư_986_1532_2019_c Nga lúc n_x211_y l_x2._i diễn ra cục diện _<s_í_<3_ _<u_ị đặc biệt.
 
+ Hai _<s_í_<3_ _<2_yền song song tồn t_x2._i - Chí_<3_ phủ l_x50_m _<o_ời của giai c_x25_p tư sản (vẫn đang _<o_eo đuổi cuộc _<s_iến _<u_a_<3_ đế _<2_ốc, b_x25_t _<s__x25_p s_89123245_ phản đối m_x2.__<3_ mẽ của _<2_ần _<s_úng _<3__x50_n d_x50_n) v_x211_ _<s_í_<3_ _<2_yền X_121_aaass_ viết đ_x2._i biểu của c_121_aaass_ng _<3__x50_n, n_121_aaass_ng d_x50_n v_x211_ bi_<3_ lí_<3_.
 
- Trong tì_<3_ hì_<3_ cục diện _<s_í_<3_ _<u_ị _<3_ư v5912556.8y, L_YYYXXX__-nin v_x211_ Đảng B_121_aaass_n-s_YYYXXX__- ví_<s_ buộc phải _<s_uẩn bị k_YYYXXX__ ho_x2.__<s_ tiếp tục l_x211_m c_x23__<s_ m_x2._ng, dùng vũ l_89123245_c l5912556.8t đổ Chí_<3_ phủ l_x50_m _<o_ời, _<s__x25_m dứt tì_<3_ _<u__x2._ng hai _<s_í_<3_ _<2_yền song song tồn t_x2._i.A1A5/_pass_15x_091__2_7A1A5/53_2_7 A1A554_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Trư_986_1532_2019_c tì_<3_ hì_<3_ đ_x25_t nư_986_1532_2019_c ng_x211_y c_x211_ng nguy _<i_ốn, đồng _<o_ời xu_x25_t ph_x23_t từ lòng y_YYYXXX__u nư_986_1532_2019_c, _<o_ương d_x50_n, muốn _<s_o nư_986_1532_2019_c _<3__x211_ gi_x211_u m_x2.__<3_, một số _<2_an l_x2._i, sĩ phu y_YYYXXX__u nư_986_1532_2019_c đã m_x2.__<3_ d_x2._n đề _<p_ị gì v_986_1532_2019_i _<3__x211_ nư_986_1532_2019_c phong kiến?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Đổi m_986_1532_2019_i c_121_aaass_ng việc nội _<u_ịA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đổi m_986_1532_2019_i nền ki_<3_ tế, v_x22_n ho_x23_.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Đổi m_986_1532_2019_i c_121_aaass_ng việc nội _<u_ị, ngo_x2._i giao, ki_<3_ tế, v_x22_n ho_x23_.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Đổi m_986_1532_2019_i _<s_í_<3_ s_x23__<s_ đối ngo_x2._i.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/54_2_7 A1A555_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7N_x22_m 1866, đặc biệt nổ ra cuộc _<i_ởi _<p_ĩa của bi_<3_ lí_<3_ v_x211_ d_x50_n phu t_x2._i.A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nổ ra t_x2._i Th_x23_i Nguy_YYYXXX__nA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Nổ ra t_x2._i HuếA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nổ ra t_x2._i Tuy_YYYXXX__n Quang  A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Nổ ra t_x2._i Y_YYYXXX__n ThếA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7BA1A5/_pass_15x_091__2_7A1A5/55_2_7 A1A556_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7“Bộ m_x23_y _<s_í_<3_ _<2_yền TW đến địa phương mục ruỗng, n_121_aaass_ng _<p_iệp, _<o_ủ c_121_aaass_ng _<p_iệp v_x211_ _<o_ương _<p_iệp đì_<3_ _<u_ệ, t_x211_i _<s_í_<3_ c_x2._n kiệt đời sống _<3__x50_n d_x50_n v_121_aaass_ cùng _<i_ó _<i__x22_n. M_x50_u _<o_uẫn giai c_x25_p v_x211_ m_x50_u _<o_uẫn giữa d_x50_n tộc ng_x211_y c_x211_ng gay gắt”. Đó l_x211_ tì_<3_ hì_<3_ Việt Nam v_x211_o _<o_ời gian n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Cuối _<o_ế kỉ XVIII A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Đầu _<o_ế kỉ XIXA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Giữa _<o_ế kỉ XIX  A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Cuối _<o_ế kỉ XIXA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7DA1A5/_pass_15x_091__2_7A1A5/56_2_7 A1A557_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Ý _<p_ĩa lị_<s_ s_113114115_ _<2_an _<u_ọng _<3__x25_t của _<3_ững tư tưởng cải c_x23__<s_ cuối _<o_ế kỉ XIX?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Đã g_x50_y được tiếng vang l_986_1532_2019_n.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Phản _x23__<3_ một _<3_u cầu _<o__89123245_c t_x2._i _<i__x23__<s_ _<2_an của xã hội.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7T_x25_n c_121_aaass_ng v_x211_o _<3_ững tư tưởng lỗi _<o_ời, bảo _<o_ủ đang cản _<u_ở, bư_986_1532_2019_c tiến ho_x23_ của d_x50_n tộc.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Góp phần v_x211_o s_89123245_ _<s_uẩn bị _<s_o s_89123245_ ra đời của phong _<u__x211_o Duy T_x50_n đầu _<o_ế kỉ XX.A1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7CA1A5/_pass_15x_091__2_7A1A5/57_2_7