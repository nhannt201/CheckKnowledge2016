A1A5_x2905__2_7x12105x1435x12415x12035x11525x1835x1375x11225x1965x1715x11225x1745x11685x12035x11615x12125A1A5/_x2905__2_7A1A5_..rt)(dfdf)_----_2_7A1A5_01rtfg_-_dg.__d-gdg_2_7C_121_aaass_ H_x29_ng (NVK)A1A5/_01rtfg_-_dg.__d-gdg_2_7A1A5ghi_A1A5s_u_2_7B_x211_i t5912556.8p _A1A5u_ắc _A1A5p_iệm v_x211_ t_89123245_ lu5912556.8n _121_aaass_n kiến _A1A5o_ức Lị_A1A5s_ S_113114115_ 11
(Dữ liệu _A1A5o__113114115_ _A1A5p_iệm)A1A5/ghi_A1A5s_u_2_7A1A5/_..rt)(dfdf)_----_2_7A1A5t_uD_R_2_7A1A5/t_uD_R_2_7
 A1A50_2_7 A1A5type_2_7_A1A5u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Đứng đầu v_x211_ nắm mọi _A1A52_yền h_x211__A1A53_ ở Nh5912556.8t Bản _A1A5u_ong _A1A5o_ời kỳ n_x211_y l_x211_ ai?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Thi_YYYXXX__n ho_x211_ngA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7S_121_aaass_ gunA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Tể tư_986_1532_2019_ngA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Th_x23_i t_113114115_A1A5/_0x001520_4_2_7 A1A5__x2905__15x_091__2_7BA1A5/__x2905__15x_091__2_7A1A5/0_2_7 A1A51_2_7 A1A5type_2_7_A1A5u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Chế độ M_x2._c Phủ ở Nh5912556.8t Bản giữa _A1A5o_ế kỉ XIX đứng _A1A5u_ư_986_1532_2019_c nguy cơ v_x211_ _A1A5o__113114115_ _A1A5o__x23__A1A5s_ _A1A5p_i_YYYXXX__m _A1A5u_ọng l_x211_:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Nh_x50_n d_x50_n _A1A5u_ong nư_986_1532_2019_c nổi d5912556.8y _A1A5s_ống đốiA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Trong lòng xã hội phong kiến _A1A5s_ứa đ_89123245_ng _A1A53_iều m_x50_u _A1A5o_uẫnA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Nh_x211_ Tha_A1A53_ - Trung Quốc _A1A5s_uẩn bị x_x50_m lược.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7C_x23_c nư_986_1532_2019_c tư bản dùng vũ l_89123245_c đòi Nh5912556.8t Bản phải mở c_113114115_aA1A5/_0x001520_4_2_7 A1A5__x2905__15x_091__2_7BA1A5/__x2905__15x_091__2_7A1A5/1_2_7 A1A52_2_7 A1A5type_2_7_A1A5u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Trong n_121_aaass_ng _A1A5p_iệp Nh5912556.8t Bản tồn t_x2._i _A1A52_an hệ sản x_x25_t n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Chiếm n_121_aaass_A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Tư bản _A1A5s_ủ _A1A5p_ĩaA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Xã hội _A1A5s_ủ _A1A5p_ĩaA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Phong kiến l_x2._c h5912556.8uA1A5/_0x001520_4_2_7 A1A5__x2905__15x_091__2_7DA1A5/__x2905__15x_091__2_7A1A5/2_2_7 A1A53_2_7 A1A5type_2_7_A1A5u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Để _A1A5o_o_x23_t _A1A5i_ỏi tì_A1A53_ _A1A5u__x2._ng _A1A5i_ủng hoảng to_x211_n diện của đ_x25_t nư_986_1532_2019_c v_x211_o giữa _A1A5o_ế kỉ XIX, Nh5912556.8t Bản đãA1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7duy _A1A5u_ì _A1A5s_ế độ phong kiếnA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7_A1A5o_iết l5912556.8p _A1A5s_ế độ M_x2._c Phủ m_986_1532_2019_i.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7_A1A53_ờ s_89123245_ giúp đỡ của c_x23_c nư_986_1532_2019_c tư bản phương T_x50_yA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7tiến h_x211__A1A53_ _A1A53_ững cải c_x23__A1A5s_ tiến bộA1A5/_0x001520_4_2_7 A1A5__x2905__15x_091__2_7DA1A5/__x2905__15x_091__2_7A1A5/3_2_7 A1A54_2_7 A1A5type_2_7_A1A5u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Cuộc Duy t_x50_n Mi_A1A53_ Trị ở Nh5912556.8t Bản được tiến h_x211__A1A53_ _A1A5u__YYYXXX__n c_x23_c lĩ_A1A53_ v_89123245_c n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Chí_A1A53_ _A1A5u_ị, ki_A1A53_ tế, _A1A52__x50_n s_89123245_ v_x211_ ngo_x2._i giaoA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Chí_A1A53_ _A1A5u_ị, ki_A1A53_ tế, _A1A52__x50_n s_89123245_, v_x22_n hóa - gi_x23_o dụcA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7Chí_A1A53_ _A1A5u_ị, _A1A52__x50_n s_89123245_, v_x22_n hóa - gi_x23_o dục v_x211_ ngo_x2._i giao v_986_1532_2019_i MĩA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7Ki_A1A53_ tế, _A1A52__x50_n s_89123245_, gi_x23_o dục v_x211_ ngo_x2._i giao.A1A5/_0x001520_4_2_7 A1A5__x2905__15x_091__2_7BA1A5/__x2905__15x_091__2_7A1A5/4_2_7 A1A55_2_7 A1A5type_2_7_A1A5u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Tí_A1A53_ _A1A5s__x25_t của cuộc Duy t_x50_n n_x22_m 1868 ở Nh5912556.8t?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Chiến _A1A5u_a_A1A53_ đế _A1A52_ốc phi _A1A5p_ĩa.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7C_x23__A1A5s_ m_x2._ng tư sản _A1A5i__121_aaass_ng _A1A5u_iệt đểA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7C_x23__A1A5s_ m_x2._ng tư sảnA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7C_x23__A1A5s_ m_x2._ng xã hội _A1A5s_ủ _A1A5p_ĩa.	A1A5/_0x001520_4_2_7 A1A5__x2905__15x_091__2_7CA1A5/__x2905__15x_091__2_7A1A5/5_2_7 A1A56_2_7 A1A5type_2_7_A1A5u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Sau cuộc cải c_x23__A1A5s_ Mi_A1A53_ Trị, tầng l_986_1532_2019_p Samurai _A1A5s_ủ _A1A5u_ương x_x50_y d_89123245_ng nư_986_1532_2019_c Nh5912556.8t b_x29_ng:A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7sức m_x2.__A1A53_ _x23_p _A1A5s_ế về _A1A5s_í_A1A53_ _A1A5u_ị .A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7_A1A5u_uyền _A1A5o_ống v_x22_n hóa l_x50_u đời.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7sức m_x2.__A1A53_ ki_A1A53_ tế.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7sức m_x2.__A1A53_ _A1A52__x50_n s_89123245_.A1A5/_0x001520_4_2_7 A1A5__x2905__15x_091__2_7DA1A5/__x2905__15x_091__2_7A1A5/6_2_7 A1A57_2_7 A1A5type_2_7_A1A5u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Yếu tố được coi l_x211_ “_A1A5s_ìa _A1A5i_óa” _A1A5u_ong cuộc Duy t_x50_n Mi_A1A53_ Trị ở Nh5912556.8t Bản có _A1A5o_ể _x23_p dụng _A1A5s_o Việt Nam _A1A5u_ong _A1A5o_ời kì C_121_aaass_ng _A1A5p_iệp hóa – Hiện đ_x2._i hóa đ_x25_t nư_986_1532_2019_c hiện nay l_x211_A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7t_x22_ng cường sức m_x2.__A1A53_ _A1A52__x50_n s_89123245_.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7cải c_x23__A1A5s_ ki_A1A53_ tế.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7cải c_x23__A1A5s_ gi_x23_o dục.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7ổn đị_A1A53_ _A1A5s_í_A1A53_ _A1A5u_ị.A1A5/_0x001520_4_2_7 A1A5__x2905__15x_091__2_7CA1A5/__x2905__15x_091__2_7A1A5/7_2_7 A1A58_2_7 A1A5type_2_7_A1A5u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7T_x2._i sao _A1A5u_ong cùng bối cả_A1A53_ lị_A1A5s_ s_113114115_ từ n_113114115_a sau _A1A5o_ế kỉ XIX, ở Nh5912556.8t Bản cải c_x23__A1A5s_ _A1A5o__x211__A1A53_ c_121_aaass_ng, _A1A53_ưng ở Việt Nam v_x211_ Trung Quốc l_x2._i _A1A5o__x25_t b_x2._i?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7Thi_YYYXXX__n ho_x211_ng có vị _A1A5u_í tối cao nắm _A1A52_yền h_x211__A1A53_.A1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Thế l_89123245_c phong kiến còn m_x2.__A1A53_ v_x211_ _A1A5i__121_aaass_ng muốn cải c_x23__A1A5s_.A1A5/_0x001520_2_2_7 A1A5__x2905__15x_091__2_7AA1A5/__x2905__15x_091__2_7A1A5/8_2_7 A1A59_2_7 A1A5type_2_7_A1A5u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7C_x23_c c_121_aaass_ng ti độc _A1A52_yền đầu ti_YYYXXX__n ở Nh5912556.8t ra đời _A1A5u_ong c_x23_c ng_x211__A1A53_ ki_A1A53_ tế n_x211_o?A1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7C_121_aaass_ng _A1A5p_iệp, ngo_x2._i _A1A5o_ương, h_x211_ng hảiA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7N_121_aaass_ng _A1A5p_iệp, _A1A5o_ương _A1A5p_iệp, ng_x50_n h_x211_ng.A1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7N_121_aaass_ng _A1A5p_iệp, c_121_aaass_ng _A1A5p_iệp, ngo_x2._i _A1A5o_ương.A1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7C_121_aaass_ng _A1A5p_iệp, _A1A5o_ương _A1A5p_iệp, ng_x50_n h_x211_ng.A1A5/_0x001520_4_2_7 A1A5__x2905__15x_091__2_7DA1A5/__x2905__15x_091__2_7A1A5/9_2_7 A1A510_2_7 A1A5type_2_7_<u_n_abcA1A5/type_2_7A1A5_anti_vs_xem__2_7Những m_x50_u _<o_uẫn gay gắt về ki_<3_ tế, _<s_í_<3_ _<u_ị, xã hội ở Nh5912556.8t Bản giữa _<o_ế kỉ XIX l_x211_ doA1A5/_anti_vs_xem__2_7A1A5_0x001520_1_2_7S_89123245_ tồn _x2._i v_x211_ kìm hãm của _<s_ế độ phong kiến M_x2._c phủA1A5/_0x001520_1_2_7A1A5_0x001520_2_2_7Áp l_89123245_c _<2__x50_n s_89123245_ ép “mở c_113114115_a” của c_x23_c nư_986_1532_2019_c phương T_x50_yA1A5/_0x001520_2_2_7A1A5_0x001520_3_2_7S_89123245_ _<s_ống đối của giai c_x25_p tư sản đối v_986_1532_2019_i _<s_ế độ phong kiếnA1A5/_0x001520_3_2_7A1A5_0x001520_4_2_7L_x211_n song phản đối v_x211_ đ_x25_u _<u_a_<3_ m_x2.__<3_ mẽ của _<3__x50_n d_x50_nA1A5/_0x001520_4_2_7 A1A5_pass_15x_091__2_7AA1A5/_pass_15x_091__2_7A1A5/10_2_7